
 /* for Linux */
 typedef signed   int32	INT;
 typedef signed   int32	SYSTIM;
 typedef signed   int32	VP_INT;
 typedef unsigned int32	UINT;
 typedef unsigned int32	UW;
 typedef unsigned int8	UB;

 /* for uITRON4.0 */

 typedef INT		ER;
 typedef INT		ID;
 typedef INT		ER_UINT;
 typedef bool		BOOL;

/*
 *  ������Хå��롼����μ����ֹ�
 */
const unsigned int SIO_ERDY_SND =   1;      /* ������ǽ������Хå� */
const unsigned int SIO_ERDY_RCV =   2;      /* �������Υ�����Хå� */

/*
 * SIGIO������������
 */
const int  LINUX_SIGIO_PRIORITY      =2;
const int  LINUX_SIGIO_STACK_SIZE =8192;


/*
 *  �ե�����ȥ���ط������
 */
const int STOP	= 23;		/* Control-S */
const int START	= 21;		/* Control-Q */

const int IXOFF_STOP	= 64;	/* buffer area size to send STOP */
const int IXOFF_START	= 128;	/* buffer area size to send START */

/*
 *  ���ꥢ�륤�󥿥ե������ɥ饤�Ф�ư�������ѤΤ�������
 *
 *  �ʲ�������ϡ��ӥå���������¤�Ȥä��Ѥ��롥
 */
const unsigned int IOCTL_NULL	=0;		/* ����ʤ� */
const unsigned int IOCTL_ECHO	=0x0001;		/* ��������ʸ���򥨥����Хå� */
const unsigned int IOCTL_CRLF	=0x0010;		/* LF �������������� CR ���ղ� */
const unsigned int IOCTL_FCSND	=0x0100;		/* �������Ф��ƥե������Ԥ� */
const unsigned int IOCTL_FCANY	=0x0200;		/* �ɤΤ褦��ʸ���Ǥ������Ƴ� */
const unsigned int IOCTL_FCRCV	=0x0400;		/* �������Ф��ƥե������Ԥ� */

/*
 *  ������μ��̤����
 *
 *  LOG_TYPE_CYC��LOG_TYPE_ASSERT �ʳ��ϡ��ǥХå��󥰥��󥿥ե�������
 *  �ͤȹ��פ��Ƥ��롥
 */
const unsigned int LOG_TYPE_INH	=	0x01;	/* ����ߥϥ�ɥ� */
const unsigned int LOG_TYPE_ISR	=	0x02;	/* ����ߥ����ӥ��롼���� */
const unsigned int LOG_TYPE_CYC	=	0x03;	/* �����ϥ�ɥ� */
const unsigned int LOG_TYPE_EXC	=	0x04;	/* CPU�㳰�ϥ�ɥ� */
const unsigned int LOG_TYPE_TEX	=	0x05;	/* �������㳰�����롼���� */
const unsigned int LOG_TYPE_TSKSTAT =	0x06;	/* �����������Ѳ� */
const unsigned int LOG_TYPE_DSP	=	0x07;	/* �ǥ����ѥå��� */
const unsigned int LOG_TYPE_SVC	=	0x08;	/* �����ӥ������� */
const unsigned int LOG_TYPE_COMMENT =	0x09;	/* ������ */
const unsigned int LOG_TYPE_ASSERT =	0x0a;	/* �����������μ��� */

const unsigned int LOG_ENTER	=	0x00;	/* ���������� */
const unsigned int LOG_LEAVE	=	0x80;	/* �и�����λ */

/*
 *  ������ν����٤����
 */
const unsigned int LOG_EMERG	=0;		/* ����åȥ�������ͤ��륨�顼 */
const unsigned int LOG_ALERT	=1;
const unsigned int LOG_CRIT	=2;
const unsigned int LOG_ERROR	=3;		/* �����ƥ२�顼 */
const unsigned int LOG_WARNING	=4;		/* �ٹ��å����� */
const unsigned int LOG_NOTICE	=5;
const unsigned int LOG_INFO	=6;
const unsigned int LOG_DEBUG	=7;		/* �ǥХå��ѥ�å����� */


const int TMAX_LOGINFO	= 6;
/* #define TMAX_LOGINFO 6 */

 const int NULL = 0;
 const int FALSE = 0;
 const int32 SERIAL_BUFSZ = 256;
 const int32 SERIAL_RCV_SEM1 = 1;
 const int32 SERIAL_SND_SEM1 = 2;
 const int32 SERIAL_RCV_SEM2 = 3;
 const int32 SERIAL_SND_SEM2 = 4;

 /*��
 	����� 
 	       factory�ǻ��ꤹ��
 	       ITRON�Ǥ���ŪAPI�ǽ�����ϥ�ɥ�˻��ꤹ��
	       �������ؿ��ǤϤʤ�

	       ������ϥ��륿���פ��Ф��ƹԤ��Τ�?
	       ����Ȥ�ġ��Υ�����Ф��ƹԤ��Τ�?

	       ʣ���Υ���ξ�硢�ġ��Υ�������ꤹ������
	       �����ͥ졼����Ϳ����ɬ�פ�����
 */


 /*
	����ߥϥ�ɥ�
		factory�ǻ��ꤹ��
		�����ߤϥ��륿���פ��Ф����������Τ�?
		������Ф����������Τ�?
				
		ʣ���Υ���ξ�硢�ġ��Υ�������ꤹ������
		�����ͥ졼����Ϳ����ɬ�פ�����
		
 	����ȥ���֥�å��ν����
		���ꥢ��ݡ��ȥ����°�����ѿ��ν�����Ǽ¸�����


 	�ݡ��Ȥν�����ϥ������³����ꤷ���Ȥ�����ޤ�

 */


 /****/

 /*
  *  ���ꥢ��ݡ��Ƚ�����֥�å�
  */

 typedef struct serial_port_initialization_block {
 	ID	rcv_semid;	/* �����Хåե������ѥ��ޥե���ID */
 	ID	snd_semid;	/* �����Хåե������ѥ��ޥե���ID */
 	char	rcv_fc_chr;	/* ����٤� START/STOP */
 } SPINIB;

/*
 *  ���ꥢ��ݡ��ȴ����֥�å������
 */
 typedef struct serial_port_control_block {
 	BOOL	openflag;	/* �����ץ�Ѥߥե饰 */
 	UINT	ioctl;		/* ư������������� */

 	UINT	rcv_read_ptr;	/* �����Хåե��ɽФ��ݥ��� */
 	UINT	rcv_write_ptr;	/* �����Хåե�����ߥݥ��� */
 	UINT	rcv_count;	/* �����Хåե����ʸ���� */
 	BOOL	rcv_stopped;	/* STOP �����ä����֤��� */

 	UINT	snd_read_ptr;	/* �����Хåե��ɽФ��ݥ��� */
 	UINT	snd_write_ptr;	/* �����Хåե�����ߥݥ��� */
 	UINT	snd_count;	/* �����Хåե����ʸ���� */
 	BOOL	snd_stopped;	/* STOP �������ä����֤��� */

 	char	rcv_buffer[SERIAL_BUFSZ];	/* �����Хåե� */
 	char	snd_buffer[SERIAL_BUFSZ];	/* �����Хåե� */
 } SPCB;

 /*
  *  ���ꥢ��I/O�ݡ��Ƚ�����֥�å�
  */
 typedef struct sio_port_initialization_block {
     UW reg_base;    /* �쥸�����Υ١������ɥ쥹 */
     UB lcr_val;     /* �⡼�ɥ쥸������������   */
     UB dlm_val;     /* �ܡ��졼�Ⱦ�̤�������   */
     UB dll_val;     /* �ܡ��졼�Ȳ��̤�������   */
     UW pinter_val;  /* ����ߵ��ĥӥå�   */    
 } SIOPINIB;

 /*
  *  ���ꥢ��I/O�ݡ��ȴ����֥�å�
  */
 typedef struct {
     VP_INT  exinf;		/* ��ĥ���� */
     BOOL    openflag;		/* �����ץ�Ѥߥե饰 */
     BOOL    sendflag;		/* ��������ߥ��͡��֥�ե饰 */
     BOOL    getready;		/* ʸ��������������� */
     BOOL    putready;		/* ʸ���������Ǥ������ */
 } SIOPCB;

 /*
  *  Linux���ߥ�졼������ѥ��ꥢ��ݡ��Ƚ�����֥�å�
  */
typedef struct serial_port_initialization_block_linux {
	ID	in_semid;	/* �����Хåե������ѥ��ޥե��� ID */
	ID	out_semid;	/* �����Хåե������ѥ��ޥե��� ID */
} SPINIBLINUX;

/*
 *  Linux���ߥ�졼������ѥ��ꥢ��ݡ��ȴ����֥�å������
 */
typedef struct serial_port_control_block_linux {
	BOOL	init_flag;	/* ������Ѥ��� */
	int	in_read_ptr;	/* �����Хåե��ɤ߽Ф��ݥ��� */
	int	in_write_ptr;	/* �����Хåե��񤭹��ߥݥ��� */
	int	out_read_ptr;	/* �����Хåե��ɤ߽Ф��ݥ��� */
	int	out_write_ptr;	/* �����Хåե��񤭹��ߥݥ��� */
	UINT	ioctl;		/* ioctl �ˤ���������� */
	BOOL	send_enabled;	/* �����򥤥͡��֥뤷�Ƥ��뤫�� */
	BOOL	ixon_stopped;	/* STOP �������ä����֤��� */
	BOOL	ixoff_stopped;	/* ���� STOP �����ä����֤��� */
	char	ixoff_send;	/* ���� START/STOP �����뤫�� */

	char	in_buffer[SERIAL_BUFSZ];	/* �����Хåե����ꥢ */
	char	out_buffer[SERIAL_BUFSZ];	/* �����Хåե����ꥢ */
} SPCBLINUX;

/* termios�ϥ��ߡ������ */
struct termios {
	int a;
};

/*
 *  Linux���ߥ�졼������ѥ��ꥢ��IO�ݡ��ȴ����֥�å������
 */
typedef struct hardware_serial_port_descripter {
	char   *path;		        /* UNIX ��ǤΥե�����̾ */
	int	   fd;		        /* �ե�����ǥ�������ץ� */
	struct termios	current_term;	/* ü��������� */
	struct termios	saved_term;    
} HWPORT;

/*
 * ����������
 */
typedef struct {
	UINT	logtype;		/* ������μ��� */
	SYSTIM	logtim;			/* ������ */
	VP_INT	loginfo[TMAX_LOGINFO];	/* ����¾�Υ����� */
} SYSLOG;


/* �������� */
signature sLogTask {
	  void main(void);	
};


/* ���������� */
signature sSysLog {
	  ER write( [in] UINT prio,  [in] SYSLOG *p_log);
	  ER_UINT read( [out] SYSLOG *p_log);
	  ER mask( [in] UINT logmask,  [in] UINT lowmask);
};



const int TCNT_SYSLOG_BUFFER = 32;


/* (�̿���)�ݡ��� */
signature sPort {
 	  ER open( void ); /* �ݡ��ȤΥ����ץ� */
 	  ER close( void ); /* �ݡ��ȤΥ����� */
 	  ER_UINT write( [in , size_is(len)] char *buf,  [in] UINT len); /* ʸ�������� */
 	  ER_UINT read( [out , size_is(len)] char *buf,  [in] UINT len); /* ʸ������� */
 	  ER ctl( [in] UINT ioctl); /* �ݡ��Ȥ����� */
};


signature sSerialPortCallBackLinux {
 	  BOOL snd( [in] VP_INT exinf);/* ���ꥢ��ݡ��Ȥ����������ǽ������Хå� */
 	  BOOL rcv( [in] VP_INT exinf); /* ���ꥢ��ݡ��Ȥ���μ������Υ�����Хå� */
};

signature sSIOPort {
 	  void open( [in] ID id , [in] VP_INT exinf);
 	  void close( [in] ID id);
 	  BOOL snd_chr( [in] char c);
 	  INT  rcv_chr( [out] char *c);
 	  void ena_cbr( [in] UINT cbrtn);
 	  void dis_cbr( [in] UINT cbrtn);
};



/* ���륿���פ���� */
[singleton] 
celltype tLogTask {
	entry sLogTask eLogTask;
	call  sSysLog cSysLog;
	call  sPort cPort;
};

[singleton] 
celltype tSysLog {
	entry sSysLog eSysLog;
	call  sPort cPort;

	  var {
	  /*
	   *  ���Ϥ��٤�������ν����١ʥӥåȥޥåס�
	    */
	    UINT	syslog_logmask;			/* ���Хåե��˵�Ͽ���٤������� */
	    UINT	syslog_lowmask;			/* ���٥���Ϥ��٤������� */
	  /*
	   *  ���Хåե��Ȥ���˥����������뤿��Υݥ���
	    */
	     SYSLOG	syslog_buffer[TCNT_SYSLOG_BUFFER];	/* ���Хåե� */
	     UINT	syslog_count;			/* ���Хåե���Υ��ο� */
	     UINT	syslog_head;			/* ��Ƭ�Υ��γ�Ǽ���� */
	     UINT	syslog_tail;			/* ���Υ��γ�Ǽ���� */
	     UINT	syslog_lost;			/* ����줿���ο� */
	  };
/*
	���ߤϡ�����ɲä���

	factory( INIT_HANDLER ,      TA_HLG, 0, tSyslog_initialize );

	
	factory( TERM_HANDLER ,      TA_HLG, 0, tSyslog_terminate );
*/
};

[singleton] 
celltype tDummySerialPort {
	entry sPort ePort;
	call  sPort cPort;
};


celltype tSerialPortLinux {
	entry sPort ePort;
	entry sSerialPortCallBackLinux eSerialPortCallBack;
	call  sSIOPort cSIOPort;

	var {
		BOOL	init_flag;	/* ������Ѥ��� */
		int	in_read_ptr;	/* �����Хåե��ɤ߽Ф��ݥ��� */
		int	in_write_ptr;	/* �����Хåե��񤭹��ߥݥ��� */
		int	out_read_ptr;	/* �����Хåե��ɤ߽Ф��ݥ��� */
		int	out_write_ptr;	/* �����Хåե��񤭹��ߥݥ��� */
		UINT	ioctl;		/* ioctl �ˤ���������� */
		BOOL	send_enabled;	/* �����򥤥͡��֥뤷�Ƥ��뤫�� */
		BOOL	ixon_stopped;	/* STOP �������ä����֤��� */
		BOOL	ixoff_stopped;	/* ���� STOP �����ä����֤��� */
		char	ixoff_send;	/* ���� START/STOP �����뤫�� */

		char	in_buffer[SERIAL_BUFSZ];	/* �����Хåե����ꥢ */
		char	out_buffer[SERIAL_BUFSZ];	/* �����Хåե����ꥢ */
	};
	attr {
		ID	in_semid;	/* �����Хåե������ѥ��ޥե��� ID */
		ID	out_semid;	/* �����Хåե������ѥ��ޥե��� ID */
	};
/* 
 �ʲ��δؿ��ϼ���ȼ����ɲä���

	 factory( INIT_HANDLER ,      TA_HLG, 0, tSerialPort_initialize );
   
*/
};

celltype tSIOPortLinux {
	entry sSIOPort eSIOPort;
	call sSerialPortCallBackLinux cSerialPortCallBack;

	var {
/* SIOPCB */
	     	VP_INT  exinf;		/* ��ĥ���� */
	     	BOOL    openflag;		/* �����ץ�Ѥߥե饰 */
	     	BOOL    sendflag;		/* ��������ߥ��͡��֥�ե饰 */
	     	BOOL    getready;		/* ʸ��������������� */
	     	BOOL    putready;		/* ʸ���������Ǥ������ */
/*	     	HWPORT    hwport;*/
		char   *path;		        /* UNIX ��ǤΥե�����̾ */
		int	   fd;		        /* �ե�����ǥ�������ץ� */
		struct termios	current_term;	/* ü��������� */
		struct termios	saved_term;    
	};

 /*
 �ʲ��δؿ��ϼ���ȼ����ɲä���

	 factory( INIT_HANDLER ,      TA_HLG, 0, tSIOPortLinux_initialize );
 	 factory( INTERRUPT_HANDLER , TA_HLG, INHNO_SIO,
 	 tSIOPortLinux_interrupt );
*/

};

/* ������Ȥ߾夲���� */

/** Log���� **/
cell tSysLog SysLog;
cell tSerialPortLinux tSerialPortLinux;

cell tLogTask LogTask {
     cSysLog = SysLog.eSysLog;
     cPort = SerialPortLinux.ePort;
};

/** DummySerialPort���� **/
cell tSerialPortLinux SerialPortLinux;

cell tDummySerialPort DummySerialPort {
     cPort = SerialPortLinux.ePort;
};

/** SysLog���� **/
cell tSysLog SysLog {
	cSIOPort = SIOPortLinux.eSIOPort;
};

/* SerialPortLinux���� */
cell tSIOPortLinux SIOPortLinux;

cell tSerialPortLinux SerialPortLinux {
	cSIOPort = SIOPortLinux.eSIOPort;

	/* var */
	init_flag = FALSE;	/* ������Ѥ��� */
	in_read_ptr = 0;	/* �����Хåե��ɤ߽Ф��ݥ��� */
	in_write_ptr = 0;	/* �����Хåե��񤭹��ߥݥ��� */
	out_read_ptr = 0;	/* �����Хåե��ɤ߽Ф��ݥ��� */
	out_write_ptr = 0;	/* �����Хåե��񤭹��ߥݥ��� */
	ioctl = 0;		/* ioctl �ˤ���������� */
	send_enabled = FALSE;	/* �����򥤥͡��֥뤷�Ƥ��뤫�� */
	ixon_stopped = FALSE;	/* STOP �������ä����֤��� */
	ixoff_stopped = FALSE;	/* ���� STOP �����ä����֤��� */
	ixoff_send = FALSE;	/* ���� START/STOP �����뤫�� */

	in_buffer = { 0 };	/* �����Хåե����ꥢ */
	out_buffer = { 0 };	/* �����Хåե����ꥢ */

	/* attr */
	in_semid = SERIAL_RCV_SEM1;
	out_semid =  SERIAL_SND_SEM1;
/*
	factory(CRE_SEM , SERIAL_RCV_SEM1, { TA_TPRI, 0, 1 });
	factory(CRE_SEM , SERIAL_SND_SEM1, { TA_TPRI, 1, 1 });
*/
};

/* SIOPortLinux���� */
/**** cell tSerialPortLinux SerialPortLinux; ****/

cell tSIOPortLinux SIOPortLinux {
	cSerialPortCallBack = SerialPortLinux.eSerialPortCallBack;

     	exinf = FALSE;		/* ��ĥ���� */
 	openflag = FALSE;		/* �����ץ�Ѥߥե饰 */
	sendflag = FALSE;		/* ��������ߥ��͡��֥�ե饰 */
	getready = FALSE;		/* ʸ��������������� */
	putready = FALSE;		/* ʸ���������Ǥ������ */

	/* attr */
/*
 	reg_base = ST16C_CHB;
	lcr_val = LCR_VAL; 
	dlm_val = DLM_VAL; 
	dll_val = DLL_VAL; 
	pinter_val = PINTER_PINT7E;
*/
/*
      siopinib = { {ST16C_CHB, LCR_VAL, DLM_VAL, DLL_VAL, PINTER_PINT7E},
 		   {ST16C_CHA, LCR_VAL, DLM_VAL, DLL_VAL, PINTER_PINT6E}
 		   };
*/
/*	
	 factory( INIT_HANDLER ,      TA_HLG, 0, SIOPortLinux_initialize );
*/

};









