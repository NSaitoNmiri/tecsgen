/*
 * $BF1$8%;%k%?%$%W$N%;%k$rD>Ns$K7k9g$9$k%1!<%9(B
 *  #647, #716, #733
 */

import_C( "tecs.h" );

signature sLinkedResource{
    void main(void);
};

[active]
celltype tOSEKResource{
    [optional]
		call sLinkedResource cLinkedResource[];  /* $BG[Ns(B */
    [optional]
		call sLinkedResource cLinkedResource2;   /* $BHsG[Ns(B */
    entry sLinkedResource eLinkedResource[];
    entry sLinkedResource eLinkedResource_2;
	attr{
		char_t *name = C_EXP( "\"$cell$\"" );
		int16_t	nest_max;
	};
	var{
		int32_t	nest;
	};
};

cell tOSEKResource OSEKResource{
    cLinkedResource[] = OSEKResource_3.eLinkedResource_2;
    cLinkedResource[] = OSEKResource_2.eLinkedResource_2;
    cLinkedResource[] = OSEKResource.eLinkedResource[0];
	nest_max = 5;
};

cell tOSEKResource OSEKResource_2{
    cLinkedResource2 = OSEKResource_2.eLinkedResource_2;
	nest_max = 3;
};

cell tOSEKResource OSEKResource_3{
    cLinkedResource2 = OSEKResource_3.eLinkedResource[1];
	nest_max = 2;
};

[singleton, active]
celltype tMain {
	call sLinkedResource cLinkedResource;
};

cell tMain Main {
	cLinkedResource = OSEKResource.eLinkedResource[0];
};
