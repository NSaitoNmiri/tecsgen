typedef int32 ER;

signature sSig1 {
  ER func1( [in]int32 arg1, [out]int32 *res );
};

signature sSig2 {
  ER func1( [in]int32 arg1, [out]int32 *res );
};

signature sSig3 {
  ER func1( [in]int32 arg1, [out]int32 *res );
};

celltype tCtR1 {
  entry sSig3 eEnt;
};

celltype tCtR2 {
  call sSig2 cCall2;
  call sSig3 cCall3;
  entry sSig1 eEnt;
};

celltype tCtOuter {
  call sSig1 cCall;
  entry sSig2 eEnt;
};

/* rRegion2 ��и��� specifier ����� */
[to_through(rRegion2, TracePlugin, ""),
out_through(TracePlugin,"")]
region rRegion2 {
  /* �ץ�ȥ�������� */
  cell tCtR2 r2cell;
};

/* rRegion1 ��и��� specifier ����� */
[in_through(TracePlugin, "")]     /* ���ιԤ������ sSig3 ���Ф��� Trace ���뤬2��ľ������� */
region rRegion1{
  /* �ץ�ȥ�������� */
  cell tCtR1 r1cell;
};

cell tCtOuter outer {
  cCall = r2cell.eEnt;
};

/* �����ʺƽи��ˤǤ� specifier �����Ǥ��ʤ� */
region rRegion1 {
  cell tCtR1 r1cell {
  };
};

/* �����ʺƽи��ˤǤ� specifier �����Ǥ��ʤ� */
region rRegion2 {
  cell tCtR2 r2cell {
   cCall2 = outer.eEnt;
   cCall3 = r1cell.eEnt;
  };

  region rRegionInner {
    cell tCtR2 r2cellInner {
      cCall2 = outer.eEnt;
      cCall3 = r1cell.eEnt;
    };
  };

};


