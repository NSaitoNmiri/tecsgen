
/* 3 => 4
 * ����������Ӵؿ��Υ�͡���
 */
import_C( "cygwin_tecs.h" );

signature sSig {
	void func( void );
	void func2( void );
	void func3( void );
};


signature sSig2 {
	void funcX( void );    // func  ==> funcX
	void funcX2( void );   // func2 ==> funcX2
	void funcX3( void );   // funcX3 ����
};

celltype tCelltype {
//	entry sSig eEnt;
	entry sSig2 eEntX;   // eEnt2 ==> eEntX
};

[active]
celltype tCelltype2 {
	call sSig2  cCall;
};

cell tCelltype Cell {
};

cell tCelltype2 Cell2 {
	cCall = Cell.eEntX;
};
