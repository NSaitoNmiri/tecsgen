import_C( "cygwin_tecs.h" );

struct tTag {
	int		a;
	int		b;
};
struct tTag2 {
	int		a;
	int		b;
};

celltype tCelltype {
	attr {
		struct tTag		sta = { 1, 2 };
		struct tTag2	sta2 = { 1, 2 };
		// int		*a			 = { 11, 12 };	// ����������ɤ��Фʤ���C����ѥ���ǥ��顼��
		int		sz			= 2;
		// int		sz;
	};
	var {
		struct tTag stv  = { 3, 4 };
		// struct tTag stv2 = sta;			// ������������ Ruby �㳰

		// int		*av = a;				// ������������ Ruby �㳰
		// int		*av2 = { 1, 2 };		// ����������ɤ��Фʤ�( C����ѥ���ǥ��顼)
		[size_is(sz)]
			int		*sz_array1;
		[size_is(sz)]
			int		*sz_array2 = { 1, 2 };	// tecsgen �������������� sz �����Ĥ��餺���顼
	};
};

cell tCelltype Cell0{
};
cell tCelltype Cell1{
	// sz = 1;     ���顼 ����������Ǥ�����¿������
};
cell tCelltype Cell2{
	sz = 2;
};
