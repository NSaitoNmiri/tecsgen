/* import_C( "tecs.h" ); */

typedef int32_t ER;
typedef int32_t TMO;

signature sAlloc {
	ER  alloc( [in]int32_t size, [out]void **p );
	ER  dealloc( [in]const void *p );
};

signature sAllocTMO {
	ER  alloc( [in]int32_t size, [out]void *p, [in]TMO tmo );
	ER  dealloc( [in]const void *p );
};

celltype tAlloc {
	entry sAlloc eA;
	attr {
		int32_t  size = 8192;
	};
	var {
		[size_is(size)]
			int8_t  *buffer;
	};
};

cell tAlloc alloc {
};

signature sSendRecv {
	/* ���δؿ�̾�� send, receive ��ȤäƤ��ޤ��� allocator ����Ǥ��ʤ� */
	ER snd( [send(sAlloc),size_is(sz)]int8_t *buf, [in]int32_t  sz );
	ER rcv( [receive(sAlloc),size_is(*sz)]int8_t **buf, [out]int32_t  *sz );
};

celltype tTestComponent {
	entry  sSendRecv eS;
	entry  sSendRecv eA[2];
};

[allocator(
	eS.snd.buf=alloc.eA,
/* 	eS.rcv.buf=alloc.eA, */
	eA[0].snd.buf=alloc.eA,
	eA[1].snd.buf=alloc.eA,
	eA[0].rcv.buf=alloc.eA/* ,
	eA[1].rcv.buf=alloc.eA */
)]
cell tTestComponent comp{
};

[singleton, active]
celltype tTestClient {
	call   sSendRecv cS;
	call   sSendRecv cA[2];
};

cell tTestClient cl {
	cS = comp.eS;
	cA[0] = comp.eA[0];
	cA[1] = comp.eA[1];
};

/**** �������������˥��㥨�顼 ****/

signature sAllocErr1 {
	ER  alloc( [in]int32_t size, [out]void *p );   // ��ťݥ���
	ER  dealloc( [in]const int p );                // �ݥ��󥿤Ǥʤ�
};

signature sSendRecvErr1 {
	/* ���δؿ�̾�� send, receive ��ȤäƤ��ޤ��� allocator ����Ǥ��ʤ� */
	ER snd( [send(sAllocErr1),size_is(sz)]int8_t *buf, [in]int32_t  sz );
	ER rcv( [receive(sAllocErr1),size_is(*sz)]int8_t **buf, [out]int32_t  *sz );
};

/**** �������������˥��㥨�顼 ****/

signature sAllocErr2 {
	ER  alloc( [in]const int32_t **size );   // out �Ǥʤ�
	ER  dealloc( [out]const int *p );   // in �Ǥʤ�
};

signature sSendRecvErr2 {
	/* ���δؿ�̾�� send, receive ��ȤäƤ��ޤ��� allocator ����Ǥ��ʤ� */
	ER snd( [send(sAllocErr2),size_is(sz)]int8_t *buf, [in]int32_t  sz );
	ER rcv( [receive(sAllocErr2),size_is(*sz)]int8_t **buf, [out]int32_t  *sz );
};

/**** �������������˥��㥨�顼 ****/

signature sAllocErr3 {
	ER  alloc( [out]int32_t ***size );   // ���ťݥ���
	ER  dealloc( [in]const int **p );   // ��ťݥ���
};

signature sSendRecvErr3 {
	/* ���δؿ�̾�� send, receive ��ȤäƤ��ޤ��� allocator ����Ǥ��ʤ� */
	ER snd( [send(sAllocErr3),size_is(sz)]int8_t *buf, [in]int32_t  sz );
	ER rcv( [receive(sAllocErr3),size_is(*sz)]int8_t **buf, [out]int32_t  *sz );
};

/**** �������������˥��㥨�顼 ****/

signature sAllocErr4 {
	ER  alloc( [in]int32_t sz, [out]int32_t ***size );   // ���ťݥ���
	ER  dealloc( [in]const int **p );   // ��ťݥ���
};

signature sSendRecvErr4 {
	/* ���δؿ�̾�� send, receive ��ȤäƤ��ޤ��� allocator ����Ǥ��ʤ� */
	ER snd( [send(sAllocErr4),size_is(sz)]int8_t *buf, [in]int32_t  sz );
	ER rcv( [receive(sAllocErr4),size_is(*sz)]int8_t **buf, [out]int32_t  *sz );
};

