[active]
celltype tAttr {
	attr {
		int	*a = { 1, 2 };
	};
	var {
		int	*b = a;			// Expression#eva_const2 ���㳰
		int	*c = ~ a;		// Expression#elements_eval_const ���㳰
		int	*d = ! a;		// Expression#elements_eval_const ���㳰
		int	*e = - a;		// Expression#elements_eval_const ���㳰
		int	*f = + a;		// Expression#elements_eval_const ���㳰
		int	*g = & a;		// Expression#elements_eval_const ���㳰
		int	*h = * a;		// Expression#elements_eval_const ���㳰
		int	*i = a + 2;		// Expression#elements_eval_const ���㳰
		int	*j = a - 2;		// Expression#elements_eval_const ���㳰
		int	*k = a * 2;		// Expression#elements_eval_const ���㳰
		int	*l = a / 2;		// Expression#elements_eval_const ���㳰
		int	*m = a % 2;		// Expression#elements_eval_const ���㳰
		int	*n = a ^ 2;		// Expression#elements_eval_const ���㳰
		int	*o = a && 2;	// Expression#elements_eval_const ���㳰
		int	*p = a | 2;		// Expression#elements_eval_const ���㳰
		int	*q = a || 2;	// Expression#elements_eval_const ���㳰
		int	*r = a > 2;		// Expression#elements_eval_const ���㳰
		int	*s = a < 2;		// Expression#elements_eval_const ���㳰
		int	*t = a >= 2;	// Expression#elements_eval_const ���㳰
		int	*u = a <= 2;	// Expression#elements_eval_const ���㳰
		int	*v = a == 2;	// Expression#elements_eval_const ���㳰
		int	*w = a != 2;	// Expression#elements_eval_const ���㳰
		int	*x = a >> 2;	// Expression#elements_eval_const ���㳰
		int	*y = a << 2;	// Expression#elements_eval_const ���㳰
	};
};

[active]
celltype tAttr2 {
	attr {
		int	*a = { 1, 2 };
	};
	var {
		int	*b = a;			// Expression#eva_const2 ���㳰
		int	*c = ~ a;		// Expression#elements_eval_const ���㳰
		int	*d = ! a;		// Expression#elements_eval_const ���㳰
		int	*e = - a;		// Expression#elements_eval_const ���㳰
		int	*f = + a;		// Expression#elements_eval_const ���㳰
		int	*g = & a;		// Expression#elements_eval_const ���㳰
		int	*h = * a;		// Expression#elements_eval_const ���㳰
		int	*i = 2 + a;		// Expression#elements_eval_const ���㳰
		int	*j = 2 - a;		// Expression#elements_eval_const ���㳰
		int	*k = 2 * a;		// Expression#elements_eval_const ���㳰
		int	*l = 2 / a;		// Expression#elements_eval_const ���㳰
		int	*m = 2 % a;		// Expression#elements_eval_const ���㳰
		int	*n = 2 ^ a;		// Expression#elements_eval_const ���㳰
		int	*o = 2 && a;	// Expression#elements_eval_const ���㳰
		int	*p = 2 | a;		// Expression#elements_eval_const ���㳰
		int	*q = 2 || a;	// Expression#elements_eval_const ���㳰
		int	*r = 2 > a;		// Expression#elements_eval_const ���㳰
		int	*s = 2 < a;		// Expression#elements_eval_const ���㳰
		int	*t = 2 >= a;	// Expression#elements_eval_const ���㳰
		int	*u = 2 <= a;	// Expression#elements_eval_const ���㳰
		int	*v = 2 == a;	// Expression#elements_eval_const ���㳰
		int	*w = 2 != a;	// Expression#elements_eval_const ���㳰
		int	*x = 2 >> a;	// Expression#elements_eval_const ���㳰
		int	*y = 2 << a;	// Expression#elements_eval_const ���㳰
	};
};


