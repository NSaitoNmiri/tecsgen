import_C( "tecs.h" );

struct tagST {
	int32_t  a;
};

signature sSig{
  void func( void );
  int32_t func2( [in]int32_t arg );
  struct tagST func3( [in]struct tagST a );
};

/*** 1.ñ�쥻���Ŭ�� ***/
// ñ�쥻���Ŭ�� (VMT ���׺�Ŭ����������ȥ����׺�Ŭ����ޤ�)
// ����¦�Υ��뤬��Ĥǡ��ݡ��Ȥ��Ĥ���

celltype tSingleCellOptimizeCaller {
	[optional]	call sSig cCall;
	[optional]	call sSig cWhite[];
	[optional]	call sSig cBlack[];
	[optional]	call sSig cBrown[];
	entry       sSig eEnt;
};

celltype tSingleCellOptimizeCallee {
	entry sSig eEnt;
};

// �Ƥ�¦���� 1����
cell tSingleCellOptimizeCallee SingleCellOptimizeCallee;

cell tSingleCellOptimizeCaller SingleCellOptimizeCaller {
//	cCall = SingleCellOptimizeCallee.eEnt;
};
// ����¦����
cell tSingleCellOptimizeCallee SingleCellOptimizeCallee {
};
// �Ƥ�¦���� 2����
cell tSingleCellOptimizeCaller SingleCellOptimizeCaller2 {
//	cCall = SingleCellOptimizeCallee.eEnt;
};

/*** 2. VMT ���׺�Ŭ�� ***/
// ����¦�Υ��뤬��Ĥ���������������

celltype tVMTUselessOptimizeCaller {
	[optional]
		call sSig cCall;
	entry sSig eEnt;
};

celltype tVMTUselessOptimizeCallee {
	entry sSig eEnt[2];
	attr {
		int32_t  attribute = 100;
	};
};

// ����¦����
cell tVMTUselessOptimizeCallee VMTUselessOptimizeCallee;

// �Ƥ�¦���� 1����
cell tVMTUselessOptimizeCaller VMTUselessOptimizeCaller {
  cCall = VMTUselessOptimizeCallee.eEnt[0];
};
// �Ƥ�¦���� 2����
cell tVMTUselessOptimizeCaller VMTUselessOptimizeCaller2 {
  cCall = VMTUselessOptimizeCallee.eEnt[1];
};
// ����¦����
cell tVMTUselessOptimizeCallee VMTUselessOptimizeCallee {
};

/*** VMT ���׺�Ŭ��&������ȥ����׺�Ŭ�� ***/
// ����¦�Υ��뤬ʣ��������ñ��Υ��륿����

celltype tSkeltonUselessOptimizeCaller {
	[optional]
		call sSig cCall;
	entry sSig eEnt;
};

celltype tSkeltonUselessOptimizeCallee {
  entry sSig eEnt;
  attr {
	  int32_t  attribute = 100;
  };
};

// ����¦����
cell tSkeltonUselessOptimizeCallee SkeltonUselessOptimizeCallee;
cell tSkeltonUselessOptimizeCallee SkeltonUselessOptimizeCallee2;

// �Ƥ�¦���� 1����
cell tSkeltonUselessOptimizeCaller SkeltonUselessOptimizeCaller {
  cCall = SkeltonUselessOptimizeCallee.eEnt;
};
// �Ƥ�¦���� 2����
cell tSkeltonUselessOptimizeCaller SkeltonUselessOptimizeCaller2 {
  cCall = SkeltonUselessOptimizeCallee2.eEnt;
};
// ����¦����
cell tSkeltonUselessOptimizeCallee SkeltonUselessOptimizeCallee {
};
cell tSkeltonUselessOptimizeCallee SkeltonUselessOptimizeCallee2 {
};

[singleton]
celltype tMain {
	call sSig cMain[];
};
/*cell tMain Main{
	cMain[] = SingleCellOptimizeCaller.eEnt;
	cMain[] = VMTUselessOptimizeCaller.eEnt;
    cMain[] = SkeltonUselessOptimizeCallee.eEnt;
    cMain[] = SkeltonUselessOptimizeCallee2.eEnt;
	};*/

celltype tCPArray {
	[optional]
		call sSig cCall[3];
	entry sSig eEnt;
};
cell tCPArray CPArray1{
};
cell tCPArray CPArray2{
	cCall[0] = SingleCellOptimizeCaller.eEnt;
	cCall[1] = VMTUselessOptimizeCaller.eEnt;
};
cell tCPArray CPArray3{
	cCall[2] = VMTUselessOptimizeCaller.eEnt;
};

celltype tNCPArray {
	[optional]
		call sSig cCall[];    // �ƤӸ��������ǿ�̤����
};
cell tNCPArray NCPArray1{
};

cell tNCPArray NCPArray2{
	cCall[] = SingleCellOptimizeCaller.eEnt;
	cCall[] = VMTUselessOptimizeCaller.eEnt;
};

[singleton]
composite tComposite {
	call sSig cMain[];
	[optional]
		call sSig cCall[3];

	cell tMain Main{
//		cMain = composite.cMain;
		cMain => composite.cMain;
	};
	cell tCPArray CPArray {
		cCall => composite.cCall;
	};
};

cell tComposite Comp
{
	cMain[] = SingleCellOptimizeCaller.eEnt;
	cMain[] = VMTUselessOptimizeCaller.eEnt;
    cMain[] = SkeltonUselessOptimizeCallee.eEnt;
    cMain[] = SkeltonUselessOptimizeCallee2.eEnt;
    cMain[] = CPArray1.eEnt;
    cMain[] = CPArray2.eEnt;
    cMain[] = CPArray3.eEnt;
};
