import_C( "cygwin_tecs.h" );

/*
 *  ���������Τ�ƤӽФ�����Υ����˥���
 */
signature sTaskBody {
	void	main(void);
};

/*
 *  �������㳰�����롼�������Τ�ƤӽФ������˥���
 */
signature sTaskExceptionBody {
	void	main([in] TEXPTN pattern);
};

[active]
celltype tTask {

          	   call	sTaskBody	cBody;  /* ���������� */
    [optional] call	sTaskExceptionBody	cExceptionBody;
									/* �������㳰�����롼�������� */
	attr{
		// ID				id = C_EXP("TSKID_$id$");
		/*
		 *  TA_NULL     0x00U   �ǥե������
		 * 	TA_ACT		0x01U	���������������˥�������ư����
		 */
		ATR		taskAttribute = C_EXP("TA_NULL");
		/*
		 * �������㳰�����롼����˻���Ǥ���°���Ϥʤ�����
		 * TA_NULL����ꤹ��
		 */
		ATR		exceptionAttribute = C_EXP("TA_NULL");
		PRI		priority;
		SIZE	stackSize;
		char_t *name = C_EXP( "\"$id$\"" );
	};
};
[context("task")]
signature sKernel{

//	ER		sleep(void);
//	ER		sleepTimeout([in] TMO timeout);
	ER		delay([in] RELTIM delay_time);

	ER		exitTask(void);
//	ER		getTaskId([out]ID *p_task_id);

//	ER		rotateReadyQueue([in] PRI task_priority);
	
	ER		getTime([out]SYSTIM *p_system_time);
	ER		getMicroTime([out]SYSUTM *p_system_micro_time);
	
//	ER		lockCpu(void);
//	ER		unlockCpu(void);
//	ER		disableDispatch(void);
//	ER		enableDispatch(void);
//	ER      disableTaskException(void);
//	ER      enableTaskException(void);
//	ER      changeInterruptPriorityMask([in] PRI interrupt_priority);
//	ER      getInterruptPriorityMask([out] PRI *p_interrupt_priority);

	ER		exitKernel(void);
//	bool_t	senseContext(void);
//	bool_t	senseLock(void);
//	bool_t	senseDispatch(void);
//	bool_t	senseDispatchPendingState(void);
//	bool_t	senseKernel(void);
};
[context("non-task")]
signature siKernel {

//	ER      getTaskId([out]ID *p_task_id);
//	ER		rotateReadyQueue([in] PRI task_priority);
	ER		getMicroTime([out]SYSUTM *p_system_micro_time);
	
//	ER      lockCpu(void);
//	ER      unlockCpu(void);

//	ER		exitKernel(void);
//	bool_t	senseContext(void);
//	bool_t	senseLock(void);
//	bool_t	senseDispatch(void);
//	bool_t	senseDispatchPendingState(void);
//	bool_t	senseKernel(void);

	/* CPU�㳰�ϥ�ɥ���ǻ��Ѥ��� */
//	bool_t	senseDispatchPendingStateCPU([in] const void * p_exception_infomation);
//	bool_t	senseTaskExceptionPendingStateCPU([in] const void * p_exception_infomation);
};

[singleton]
celltype tKernel{
	[inline] entry sKernel  eKernel;
	[inline] entry siKernel eiKernel;
};
/*
 * ���ޥե��Υ����˥���ʥ���������ƥ������ѡ�
 */
signature sSemaphore{
	ER 		signal(void);
	ER 		wait(void);
	ER 		waitPolling(void);
	ER 		waitTimeout([in] TMO timeout);
	ER 		initialize(void);
	ER 		refer([out] T_RSEM *pk_semaphore_status);
};

/*
 *  ���ޥե��Υ����˥�����󥿥�������ƥ������ѡ�
 */
[context("non-task")]
signature siSemaphore {
	ER 		signal(void);
};
/*
 * ���ޥե��Υ��륿�������
 */
celltype tSemaphore{
	[inline]entry  sSemaphore   eSemaphore; /* ���ޥե����ʥ���������ƥ������ѡ�*/
	[inline]entry  siSemaphore  eiSemaphore;/* ���ޥե������󥿥�������ƥ������ѡ�*/
	
	attr {
		ID      id = 0/* = C_EXP( "SEMID_$id$" )*/;
		[omit]  ATR attribute;
		[omit]  uint32_t count;
		[omit]  uint32_t max =1;

	};
	var {
		pthread_mutex_t  mutex = C_EXP( "PTHREAD_MUTEX_INITIALIZER" );
	};

//	factory {
//		write( "tecsgen.cfg", "CRE_SEM(%s, { %s, %s, %s });", id, attribute, count, max);
//	};
//	FACTORY{
//		write( "$ct$_factory.h","#include \"kernel_cfg.h\"" );
//	};
};

/*
 *  ���٥�ȥե饰�Υ����˥���ʥ���������ƥ������ѡ�
 */
signature sEventflag{
	ER set([in] FLGPTN set_pattern);
	ER clear([in] FLGPTN clear_pattern);
	ER wait([in] FLGPTN wait_pattern, [in] MODE wait_flag_mode, [out] FLGPTN *p_flag_pattern);
	ER waitPolling([in] FLGPTN wait_pattern, [in] MODE wait_flag_mode, [out] FLGPTN *p_flag_pattern);
	ER waitTimeout([in] FLGPTN wait_pattern, [in] MODE wait_flag_mode, [out] FLGPTN *p_flag_pattern, [in] TMO timeout);

	ER initialize(void);
	ER refer([out]T_RFLG *pk_eventflag_status);
};
/*
 *  ���٥�ȥե饰�Υ����˥�����󥿥�������ƥ������ѡ�
 */
[context("non-task")]
signature siEventflag {
	ER set([in] FLGPTN set_pattern);
};
/*
 *  ���٥�ȥե饰
 */
celltype tEventflag{
	/*[inline]*/ entry  sEventflag   eEventflag; /* ���٥�ȥե饰���ʥ���������ƥ������ѡ�*/
	/*[inline]*/ entry  siEventflag  eiEventflag;/* ���٥�ȥե饰�����󥿥�������ƥ������ѡ�*/
	
	attr {
		ID      id = 0 /*C_EXP( "FLGID_$id$" )*/;
		/*
		 * TA_NULL �ǥե�����͡�FIFO�Ԥ���
         * TA_TPRI �Ԥ�����򥿥�����ͥ���ٽ�ˤ���
         * TA_WMUL ʣ���Υ��������ԤĤΤ����
         * TA_CLR  ���������Ԥ�������˥��٥�ȥե饰�򥯥ꥢ����
		 */
		[omit]  ATR attribute = C_EXP("TA_NULL");
		/*
		 * ���٥�ȥե饰�Υӥåȥѥ�����ν����
		 */
		[omit]  FLGPTN flagPattern;
	};
	var {
		pthread_mutex_t   mutex      = C_EXP( "PTHREAD_MUTEX_INITIALIZER" );
//		pthread_mutex_t   cond_mutex = C_EXP( "PTHREAD_MUTEX_INITIALIZER" );
		pthread_cond_t    cond       = C_EXP( "PTHREAD_COND_INITIALIZER" );
		pthread_once_t    once       = C_EXP( "PTHREAD_ONCE_INIT" );
		FLGPTN            pattern    = flagPattern;
	};

//	factory {
//		write( "tecsgen.cfg", "CRE_FLG(%s, { %s, %s});", id, attribute, flag_pattern);
//	};
//	FACTORY{
//		write( "$ct$_factory.h", "#include \"kernel_cfg.h\"" );
//	};
};


/*
 *  �ǡ������塼�����뤿��Υ����˥���ʥ���������ƥ������ѡ�
 */
signature sDataqueue {
	/*�ǡ������塼������*/
	ER 		send([in] intptr_t data);
	ER 		sendPolling([in] intptr_t data);
	ER 		sendTimeout([in] intptr_t data, [in]TMO timeout);
	ER 		sendForce([in] intptr_t data);
	/*�ǡ������塼�μ���*/
	ER 		receive([out] intptr_t *p_data);
	ER 		receivePolling([out] intptr_t *p_data);
	ER 		receiveTimeout([out] intptr_t *p_data, [in]TMO timeout);
	
	ER 		initialize(void);
	ER 		refer([out] T_RDTQ *pk_dataqueue_status);
};
/*
 *  �ǡ������塼�����뤿��Υ����˥�����󥿥�������ƥ������ѡ�
 */
[context("non-task")]
signature siDataqueue {
	ER 		sendPolling([in] intptr_t data); 
	ER 		sendForce([in] intptr_t data);
};
/*
 *  �ǡ������塼
 */
celltype tDataqueuePeer {
	[inline] entry  sDataqueue   eDataqueue; /* �ǡ������塼���ʥ���������ƥ������ѡ�*/
	[inline] entry  siDataqueue  eiDataqueue;/* �ǡ������塼�����󥿥�������ƥ������ѡ�*/
	call  sSemaphore  cInitializing;
	
	attr {
//		ID      id = C_EXP( "DTQID_$id$" );
		/*
		 * TA_NULL �ǥե�����͡�FIFO���
		 * TA_TPRI �����Ԥ�����򥿥�����ͥ���ٽ�ˤ���
		 */
		ATR     attribute = C_EXP( "TA_NULL" );
		uint_t  count = 1;
		void    *pdqmb = C_EXP( "NULL" );
	};
	var {
		int_t   fd[2];   // pipe �Υǥ�������ץ��ֹ�
		bool_t  b_init;
	};

};

composite tDataqueue {
	entry  sDataqueue   eDataqueue; /* �ǡ������塼���ʥ���������ƥ������ѡ�*/
	entry  siDataqueue  eiDataqueue;/* �ǡ������塼�����󥿥�������ƥ������ѡ�*/
	attr {
		uint_t	count;
	};

	cell tSemaphore Semaphore {
		count = 1;
		max = 1;
		attribute = C_EXP("TA_NULL");
	};
	cell tDataqueuePeer Peer {
		cInitializing = Semaphore.eSemaphore;
		count = composite.count;
	};
	composite.eDataqueue  => Peer.eDataqueue;
	composite.eiDataqueue => Peer.eiDataqueue;
};
