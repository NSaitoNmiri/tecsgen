/*
 * ����ե��������Υƥ���
 */

import_C( "cygwin_tecs.h" );
import( "cygwin_kernel.cdl" );

signature sAlloc {
	ER  alloc( [in]int32_t sz, [out]void **p );
	ER  dealloc( [in]const void *p );
};

signature sSig {
	ER  func( [send(sAlloc)]int32_t *a );
	ER  func2( [send(sAlloc),size_is(sz)]int8_t *buf, [in]int32_t sz );
};

celltype tAlloc {
	entry sAlloc eA;
	attr {
		int32_t  num;
	};
};

celltype tCt1 {
	entry sSig eEnt;
	attr {
		int32_t  num;
	};
};

[active,singleton]
celltype tCt2 {
	call sSig cCall[];
};

// composite ��Υ���ե�������
composite tCompAlloc {

	entry sAlloc eAlloc;
	[allocator(
		func.a=eAlloc,
		func2.buf=eAlloc)]
	entry sSig  eEntExt;
	attr {
		int32_t  num;
	};

	[allocator(
		eEnt.func.a=Alloc.eA,
		eEnt.func2.buf=Alloc.eA)]
	cell tCt1 Cell1 {
		num = composite.num;
	};

	cell tAlloc Alloc{
		num = composite.num;
	};

	cell tAlloc Alloc2{
		num = composite.num;
	};

	composite.eEntExt => Cell1.eEnt;
	composite.eAlloc  => Alloc.eA;
	// composite.eAlloc  => Alloc2.eA;
};


// --------  2���� -------

cell tCt2 Cell2{
	cCall[] = CompAlloc.eEntExt;
	cCall[] = CompAlloc2.eEntExt;
};

cell tCompAlloc CompAlloc{
	num = 1;
};

cell tCompAlloc CompAlloc2{
	num = 2;
};

// ����ե��������κƵ�Ū composite ��
//**********
composite tCompAllocSuper {
	[allocator(func.a=eAlloc,
			   func2.buf=eAlloc)]
	entry	sSig	eEntExt2;
	entry	sAlloc	eAlloc;
	attr {
		int32_t  num;
	};	
	
	cell tCompAlloc CellIn{
		num = composite.num;
	};
	cell tAlloc Alloc{
		num = composite.num;
	};
	composite.eEntExt2 => CellIn.eEntExt;
	composite.eAlloc   => CellIn.eAlloc;
	// composite.eAlloc   => Alloc.eA;
};

cell tCompAllocSuper CompAllocSuper{
	num = 10;
};

[active,singleton]
celltype tCt3 {
	call sSig cCall;
};

cell tCt3 Cell3{
	cCall = CompAllocSuper.eEntExt2;
};

// **********/

/*****

����������������

���������� composite ����¦���֤��������send/receive �����Υ����������礵������������������������

���͡�
�����������μ������ϳ����������ʤ��ƤϤʤ�ʤ�
��composite �μ�����������ǡ����������λ����Ԥ�

��ͳ��
�����󥿥ե��������򸫤������ǡ�������礵��Ƥ��뤳�Ȥ��狼��
���Ƶ�Ū�� composite ��Ʊ����ˡ�Ǽ¸��Ǥ���

������
tCompAlloc ��������줿�Ȥ�
��tCompAlloc �� new_port �ˤ�����
  ���⤷��(3) �ˤ�����������������(2) �����ꤵ��Ƥ���ʤ��
    ��(3�ˤΥ����å��ˤ�����
        (2)�κ��դΰ����� (3) �Υ����˥����¸�ߤ���
        (2)�α���eAlloc �� signature �� func.a �� send �� alloc �Ȱ��פ��뤳�Ȥ�����å�
        @internal_allocator_list �����
��tCompAlloc �� new_join �ˤ�����
  ���⤷����3�ˤ� func.a �˥�졼��������/����������������ʤ���С��������������ؤ� new_join ��Ԥ�
��tCompAlloc �� end_of_parse �ˤ�����
  (2) �Υ������������ (5) ������������������̷�⤬�ʤ����Ȥγ�ǧ
  ��(3) �ˤĤ���
    (2) �α��� eAlloc �� (1) �� (9) �Ȥ��ɤ������η���� Alloc.eAlloc ������
    (3) �� (8) �� (6) �Ȥ��ɤ����� Cell1 ��õ��
    ���⤷ Cell1 �� alloc_list �����Ƥ� eEnt_func_a ������С�
        Alloc.eAlloc �˰��פ��뤳�Ȥ��ǧ����
    ���ʤ���Х��顼

tCompAlloc �Υ��뤬�������줿�Ȥ�
��Cell#expand �ˤ�
  ��alloc_list �ˡ�get_allocator_list �˴�Ť��ơ� (2) �η���ä���

@internal_allocator_list ���ѹ�
   @internal_allocator_list ����������ؤη��ˤʤäƤ���������������˲����
   ���������ľ�ܷ�礹��褦�� alloc_list ����������Ƥ�������composite �Υ���Υ��������μ������ؤΤ�Τ��ѹ�
   ��CompositeCelltype#new_join ���� CompositeCelltype#new_port �ذܤ�
   ��Cell#expand

�����ε�Ͽ
��bnf.y.rb :  composite_celltype_statement_specifier �ˤ����� alloc_list => alloc_list2
��Port#set_allocator_instance
     �������������λ���򥨥顼(S1081)�Ȥ��ʤ�

*****/

/****

composite tCompAlloc {

	[allocator(
		func.a=eAlloc,                  �� (2)
		func2.buf=eAlloc)]
	entry sSig    eEntExt;              �� (3)

	entry sAlloc  eAlloc;            �� �� (1)           // �������Ȳ�ǽ

	attr {
		int32_t  num;                   �� (4)
	};

    [allocator(                         �� (5)
		eEnt.func.a=Alloc.eAlloc,
		eEnt.func2.buf=Alloc.eAlloc)]
	cell tCt1 Cell1 {                   �� (6)
		num = composite.num;
	};

	cell tAlloc Alloc{
		num = composite.num;            �� (7)
	};

	composite.eEntExt => Cell1.eEnt;    �� (8)
	composite.eAlloc  => Alloc.eAlloc;  �� (9)
};

composite tCompAllocSuper {
	entry sAlloc  eAlloc;
	[allocator(
		func.a    = eAlloc,
		func2.buf = eAlloc)]
	entry sSig    eEntExt2;
	attr {
		int32_t  num;
	};	
	cell tCompAllocNew CellIn{
		num = composite.num;
	};
	composite.eEntExt2 => CellIn.eEntExt;
	composite.eAlloc   => CellIn..eAlloc;
};

// *****/

/****

�ڥ�졼����������

tCompRelayAlloc �� end_of_parse �ˤ�
��IF (2)����Relay ���������������ġ�
��THEN
  ��(1)  �α��դ� cCall.func.a �����뤳�Ȥ�Ĵ�٤� (signature �ΰ��פ�Ĵ�٤�)
      ���դ⤢�뤳�Ȥ�Ĵ�٤�
  ��(2) eEntExt.func.a 
     => (6) Relay.eEnt.func.a     ������б����� relay allocator ������         (a)
     => (5) Relay.cCall.func.a    ���θƤӸ��η���褬�����Ǥ��뤳�Ȥ��ǧ����  (b)
     �� (4) cCallExt.func.a

  (b) �ˤ����ơ��Ƥ� relay allocator �Ǥ����礬�����¿�ʥ�졼����
      ���ξ�� (b) �� (a) ��ή��򷫤��֤�

tCompRelayAlloc �Υ��뤬�������줿�Ȥ�
��create_relay_allocaotr �ˤ����� alloc_list ����������

composite tCompRelayAlloc {
	[allocator(	func.a    <= cCallExt.func.a,  �� (1)
				func2.buf <= cCallExt.func2.buf)]
		entry	sSig	eEntExt;               �� (2)
	call		sSig	cCallExt;              �� (3)

	cell tRelayCell Relay {                    �� (4)
		cCall => composite.cCallExt;           �� (5)
	};
	composite.eEntExt => Relay.eEnt;           �� (6)
};

// ****/
