/*
 *  TECS Generator
 *      Generator for TOPPERS Embedded Component System
 *  
 *   Copyright (C) 2008-2013 by TOPPERS Project
 *--
 *   �嵭����Ԥϡ��ʲ���(1)(4)�ξ������������˸¤ꡤ�ܥ��եȥ���
 *   �����ܥ��եȥ���������Ѥ�����Τ�ޤࡥ�ʲ�Ʊ���ˤ���ѡ�ʣ������
 *   �ѡ������ۡʰʲ������ѤȸƤ֡ˤ��뤳�Ȥ�̵���ǵ������롥
 *   (1) �ܥ��եȥ������򥽡��������ɤη������Ѥ�����ˤϡ��嵭������
 *       ��ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ��꤬�����Τޤޤη��ǥ���
 *       ����������˴ޤޤ�Ƥ��뤳�ȡ�
 *   (2) �ܥ��եȥ������򡤥饤�֥������ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ�����Ǻ����ۤ�����ˤϡ������ۤ�ȼ���ɥ�����ȡ�����
 *       �ԥޥ˥奢��ʤɡˤˡ��嵭�����ɽ�����������Ѿ�浪��Ӳ���
 *       ��̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *   (3) �ܥ��եȥ������򡤵�����Ȥ߹���ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ��ʤ����Ǻ����ۤ�����ˤϡ����Τ����줫�ξ�����������
 *       �ȡ�
 *     (a) �����ۤ�ȼ���ɥ�����ȡ����Ѽԥޥ˥奢��ʤɡˤˡ��嵭����
 *         �ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *     (b) �����ۤη��֤��̤�������ˡ�ˤ�äơ�TOPPERS�ץ������Ȥ�
 *         ��𤹤뤳�ȡ�
 *   (4) �ܥ��եȥ����������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������뤤���ʤ�»
 *       ������⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ����դ��뤳�ȡ�
 *       �ޤ����ܥ��եȥ������Υ桼���ޤ��ϥ���ɥ桼������Τ����ʤ���
 *       ͳ�˴�Ť����ᤫ��⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ�
 *       ���դ��뤳�ȡ�
 *  
 *   �ܥ��եȥ������ϡ�̵�ݾڤ��󶡤���Ƥ����ΤǤ��롥�嵭����Ԥ�
 *   ���TOPPERS�ץ������Ȥϡ��ܥ��եȥ������˴ؤ��ơ�����λ�����Ū
 *   ���Ф���Ŭ������ޤ�ơ������ʤ��ݾڤ�Ԥ�ʤ����ޤ����ܥ��եȥ���
 *   �������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������������ʤ�»���˴ؤ��Ƥ⡤��
 *   ����Ǥ�����ʤ���
 *  
 *   $Id: $
 */

import_C( "netinet/in.h" );

const	uint16_t	TINETIPV4_DEFAULT_PORT_NO  = 8931;

signature sTINETClientOpenerIPV4 {
	ER		open( [in]const T_IPV4EP *clientAddr, [in]TMO tmo );
	ER		close( [in]TMO tmo );
};

signature sIPV4AcceptCheck {
	bool_t	check( [in]const T_IPV4EP *clientAddr );
};

celltype tTINETClient {
	entry	sChannel				eC0;
	entry	sTINETClientOpenerIPV4	eOpener;
	attr {
		ID				cep_id = C_EXP( "$id$_CEPID" );
		[omit]
			uint16_t	recv_buf_size = C_EXP( "TCP_MSS" );
		[omit]
			uint16_t	send_buf_size = C_EXP( "TCP_MSS" );
	};
	FACTORY {
		write( "$ct$_factory.h", "#include \"netinet/tcp.h\"\n" );
		write( "$ct$_tecsgen.h", "#include \"tinet_cfg.h\"\n" );
		write( "tinet_tecsgen.cfg", "#include \"$ct$_factory.h\"\n" );
	};
	factory {
		write( "$ct$_factory.h", "int8_t $id$_recv_buf[%s];\n", recv_buf_size );
		write( "$ct$_factory.h", "int8_t $id$_send_buf[%s];\n", send_buf_size );
		write( "tinet_tecsgen.cfg", "TCP_CRE_CEP ($id$_CEPID, {\n"
								"	0,\n"
								"	$id$_send_buf,\n"
								"	%s,\n"
								"	$id$_recv_buf,\n"
								"	%s,\n"
								"	NULL \n"
								"	} );\n",
			   send_buf_size, recv_buf_size );
	};
};

celltype tTINETServer {

	entry	sChannel				eC1;
	entry	sServerChannelOpener	eOpener;
	[optional]
		call  sIPV4AcceptCheck  cCheck;
	attr {
		ID				cep_id = C_EXP( "$id$_CEPID" );
		ID				rep_id = C_EXP( "$id$_REPID" );
		[omit]
			int16_t		portNo  = TINETIPV4_DEFAULT_PORT_NO;
		[omit]
			uint16_t	recv_buf_size = C_EXP( "TCP_MSS" );
		[omit]
			uint16_t	send_buf_size = C_EXP( "TCP_MSS" );
	};
	FACTORY {
		write( "$ct$_factory.h", "#include \"netinet/tcp.h\"\n" );
		write( "$ct$_tecsgen.h", "#include \"tinet_cfg.h\"\n" );
		write( "tinet_tecsgen.cfg", "#include \"$ct$_factory.h\"\n" );
	};
	factory {
		write( "$ct$_factory.h", "int8_t $id$_recv_buf[%s];\n", recv_buf_size );
		write( "$ct$_factory.h", "int8_t $id$_send_buf[%s];\n", send_buf_size );
		write( "tinet_tecsgen.cfg", "TCP_CRE_REP ($id$_REPID,	{ 0, { IPV4_ADDRANY, %s } } );\n", portNo );
		write( "tinet_tecsgen.cfg", "TCP_CRE_CEP ($id$_CEPID, {0, $id$_send_buf, %s, $id$_recv_buf, %s, NULL } );\n",
				   send_buf_size, recv_buf_size );
	};
};
