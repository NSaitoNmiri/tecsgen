typedef int32_t ER;

signature sOneway {
	[oneway]
		ER  func1( [in]int32_t     inval );    /* ���� */
	[oneway]
		ER  func2( [inout]int32_t  *ioval );   /* ERROR (inout ������) */
	[oneway]
		ER  func3( [out]int32_t    *outval );  /* ERROR (out ������) */
	[oneway]
		int32_t  func4( void );                /* ERROR (ER �Ǥʤ� return ������) */
};

