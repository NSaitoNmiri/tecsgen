/*
 * ��졼���������Υƥ���
 */

import_C( "tecs.h" );

/* typedef int32_t ER;
typedef int32_t TMO; */

signature sAlloc {
	ER	alloc( [in]int32_t size, [out]void **p );
	ER	dealloc( [in]const void *p );
};

signature sAllocTMO {
	ER	alloc( [in]int32_t size, [out]void *p, [in]TMO tmo );
	ER	dealloc( [in]const void *p );
};

celltype tAlloc {
	entry sAlloc eA;
	attr {
		int32_t  size = 8192;
	};
	var {
		[size_is(size)]
			int8_t	*buffer;
		int32_t	n_alloc;
		int32_t	n_dealloc;
	};
};

cell tAlloc Alloc {
};

signature sSendRecv {
	/* ���δؿ�̾�� send, receive ��ȤäƤ��ޤ��� allocator ����Ǥ��ʤ� */
	ER	snd( [send(sAlloc),size_is(sz)]int8_t *buf, [in]int32_t  sz );
	ER	rcv( [receive(sAlloc),size_is(*sz)]int8_t **buf, [out]int32_t  *sz );
};

/*
 * ��졼��������������
 */
celltype tRelayComponent {
	/* [allocator(
	   snd.buf <= cSR.snd.buf
	   )] */   /* ����������Υ�졼����������̤���ݡ��� */
	entry  sSendRecv eA[2];

	// ��졼���������λ���
	[allocator(
			   snd.buf <= cSR.snd.buf,  /* �������Ȳ�ǽ */
			   rcv.buf <= cSR.rcv.buf
			   )]
		entry  sSendRecv eS;
	call   sSendRecv cSR;

	attr {
		char_t	*name = C_EXP( "\"$id$\"" );
	};
};

celltype tTargetComponent {
	entry	sSendRecv eS;
};

[allocator(
		   eS.snd.buf=Alloc.eA,
		   eS.rcv.buf=Alloc.eA
)]
cell tTargetComponent TargetCell {
};

[allocator(
		   // eS.snd.buf=Alloc.eA,  // ��졼���������ǻ��ꤵ���
		   // eS.rcv.buf=Alloc.eA,  // ������ͭ���ˤ���ȡ���ʣ���顼�ˤʤ�
		   eA[0].snd.buf=Alloc.eA,
		   eA[1].snd.buf=Alloc.eA,
		   eA[0].rcv.buf=Alloc.eA,
		   eA[1].rcv.buf=Alloc.eA
		   )]
cell tRelayComponent RelayCell{
	cSR = TargetCell.eS;
};

[allocator(
		   // eS.snd.buf=Alloc.eA,  // ��졼���������ǻ��ꤵ���
		   // eS.rcv.buf=Alloc.eA,  // ������ͭ���ˤ���ȡ���ʣ���顼�ˤʤ�
		   eA[0].snd.buf=Alloc.eA,
		   eA[1].snd.buf=Alloc.eA,
		   eA[0].rcv.buf=Alloc.eA,
		   eA[1].rcv.buf=Alloc.eA
		   )]
cell tRelayComponent RelayCell2{
	cSR = RelayCell.eS;
};


[singleton]
celltype tTestClient {
	call   sSendRecv cS;
	call   sSendRecv cA[2];
};

cell tTestClient Client {
	cS    = RelayCell2.eS;
	cA[0] = RelayCell.eA[0];
	cA[1] = RelayCell.eA[1];
};

[singleton]
celltype tTestOptional {
	[optional]
		call   sSendRecv cS;
};

cell tTestOptional TestOptional {};
