typedef   bool BOOL;
const bool true  = 1;  /* ̯�ʽ���� */
const bool false = 1;

celltype tBool {
  attr {
    BOOL  v  = 0;
    BOOL  v2 = {1};     /* ��̣Ū���顼�ˤʤ�ʤ������������顼�� */
  };
};

cell tBool b {
};

/*
 * NULL ��Ÿ������Ƥ��ޤ�
 * #define NULL ((const int)0)     const ������, NULL ������եꥯ��
 */
