
/* typedef int32_t ER; */

signature sMain {
	void  main(void);
};

signature sSig1 {
	ER func1( [in]int32_t arg1, [out]int32_t *res );
};

signature sSig2 {
	ER func1( [in]int32_t arg1, [out]int32_t *res );
};

signature sSig3 {
	ER func1( [in]int32_t arg1, [out]int32_t *res );
};

celltype tCtR1 {
	entry sSig3 eEnt;
};

celltype tCtR2 {
	call sSig2 cCall2;
	call sSig3 cCall3;
	entry sSig1 eEnt;
};

celltype tCtOuter {
	call    sSig1  cCall;
	entry   sSig2  eEnt;
	entry   sMain  eMain;
};

/* rRegion2 ��и��� specifier ����� */
[to_through(rRegion1),
//[to_through(rRegion1, TracePlugin, "cellEntry=\"r1cell.eEnt2 , r1cell.eEnt\""),
//[to_through(rRegion1, TracePlugin, "cellEntry=\"r1cell.eEnt2\",cellEntry=\"r1cell.eEnt\""),
//[to_through(rRegion1, TracePlugin, "cellEntry=\"r1cell.eEnt2\""),
out_through(/*TracePlugin,""*/),
in_through()]
region rRegion2 {
	/* �ץ�ȥ�������� */
	cell tCtR2 r2cell;

	// TracePlugin �ǻȤ���
	cell tSysLog  SysLogn2{
	};
	cell tKernel  Kernel{
	};
};

/* rRegion1 ��и��� specifier ����� */
region rRegion1{
	/* �ץ�ȥ�������� */
	cell tCtR1 r1cell;

	// TracePlugin �ǻȤ���
//	cell tSysLog  SysLogn1{
//	};
};

cell tCtOuter outer {
	cCall = rRegion2::r2cell.eEnt;
};

/* �����ʺƽи��ˤǤ� specifier �����Ǥ��ʤ� */
region rRegion1 {
	cell tCtR1 r1cell {
	};
};

/* �����ʺƽи��ˤǤ� specifier �����Ǥ��ʤ� */
region rRegion2 {
	cell tCtR2 r2cell {
		cCall2 = outer.eEnt;
		cCall3 = rRegion1::r1cell.eEnt;
	};

	[out_through(Plugin2,"")]
	region rRegionInner {
		cell tCtR2 r2cellInner {
			cCall2 = outer.eEnt;
			/* #327 �ƤӸ��� through �� region �� through �������˽Ф뤳�ȤΥƥ��� */
			[through(Plugin1, "" )]
				cCall3 = rRegion1::r1cell.eEnt;
		};
	};
};

[singleton,active]
celltype tMain {
	call sMain cMain;
};

cell tMain Main{
	cMain = outer.eMain;
};

