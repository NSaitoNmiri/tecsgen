
/*
 * 1. tecs_bool���Υ�����ѿ��˽���ͤ����ꤷ�ʤ���硢CB�ν�����Ҥ�{}�Ƚ��Ϥ����(��:gen/tSerialPort_tecsge.c) 
 *
 *   var �ν����̤����ν��ϥ����ɤθ��
 *
 * 2. char��������Ǥ��륻����ѿ��˽���ͤ����ꤷ�ʤ���硢CB�ν�����Ҥ�{}�Ƚ��Ϥ����(��:gen/tSerialPort_tecsge.c) 
 *
 *   ����ǤϤʤ��ݥ��󥿡�
 *   ����� var �ν����̤����ν��ϥ����ɤθ��
 *
 * 3. ��¤�Τ�����򥻥���ѿ��ˤ��ơ�����ͤ����ꤷ�ʤ���硢CB�ν�����Ҥ�{}�Ƚ��Ϥ����(��:gen/tSyslog_tecsge.c) 
 *
 *   ������Զ�硩
 *
 * 4. ���顼��å������δְ㤤(��)�����������ѤΥ���������¸�ߤ��Ƥ⡢�����������Τ�¸�ߤ��ʤ���硢��refereced but defined�פȤ������顼��å�������ɽ������롣�ʤ��ι��*.cdl����Ͽ���Ƥ��ޤ���� 
 *
 *    "reference undefined cell" ���ѹ�
 *
 * 5. ��¤�Τη�����ǡ����Ф�������������ǿ���const�ѿ��ǻ���)���Ƥ⡢global_tecsgen.h�ˤ�����ǤϤʤ���ñ����ѿ��Ȥ��ƽ��Ϥ����(��:gen/global_tecsgen.h) 
 *
 *    �����Τʤ���¤�Τ� typedef �Υ��Фν��ϥ����ɤθ��
 *    ��¤�Υ����������� struct �� typedef ��������줿���Ȥˤʤ뤬���ʤ����� typedef �Τ�������줿���Ȥˤʤ�
 *    ���Ԥ� generate.rb �� StructType �� gen_gh �ǽ��Ϥ����
 *    ��Ԥ� types.rb �� get_type_str, get_type_str_post �ˤ����Ϥ����ʤ����餬�б��Ǥ��Ƥ��ʤ��ä���
 *
 * 6. ���󥰥�ȥ�Ǥʤ������°�����ѿ���ɽ���ޥ����;ʬ��&���դ��Ƥ���(IDX���ݥ��󥿤ξ���(��:gen/tSerialPort_tecsgen.h) 
 *
 *    ���ͤȻפ��ޤ�
 *    2006.8.17 �Υߡ��ƥ��󥰤� attribute �Υ��������ޥ����ݥ��󥿤��֤��褦�ˤʤ�ޤ���
 *    http://www.toppers.jp/MEMBERS/wiki/com-wg/?2006%C7%AF8%B7%EE17%C6%FC%A5%DF%A1%BC%A5%C6%A5%A3%A5%F3%A5%B0
 *
 * 7. ���󥰥�ȥ�Ǥʤ������°�����ѿ���ɽ���ޥ������Ϥ���ʤ� 
 *
 *    ���󥰥�ȥ󥻥�ξ�硩
 *    °�����ѿ��Ͻ��Ϥ���Ƥ��ޤ���
 *    ��Ŧ���ब�狼��ޤ���Ǥ�����
 *
 * 8. signature��signed char���������Ƥ⡢�����ͥ졼����tecs_char(��󥿥����unsigned char��typdef����Ƥ���ˤ���Ϥ��롣tecs_schar(��󥿥����signed char��typdef����Ƥ���ˤ���Ϥ����ߤ�����
 *
 *    �������ΰ����ˤĤ��ơ��⤦��������ľ���Ƥ�����ꤷ�����Ǥ�
 *
 */

const int32_t TMAX_LOGINFO = 10;

typedef struct tag_syslog_t  {
	int32_t	logtype;		/* ������μ��� */
	int32_t	logtim;			/* ������ */
	int32_t	loginfo[TMAX_LOGINFO];	/* ����¾�Υ����� */  /* Bug 5 */
} syslog_t;

celltype tBugTest {
  attr {
    bool_t a = false;
    char_t *path1 = "A";
    syslog_t  sys1[ 1 ] = { {  0  }}; 	/* Bug 3 */
  };
  var {
    bool_t b;			/* Bug 1 */
    char_t *path2;		/* Bug 2 */
    syslog_t  sys2[ 2 ];	/* Bug 3 */
  };
};

cell tBugTest boolTest {
  
};

[singleton]
celltype tSingle {
  attr {
    int32_t a = 0;
  };
  var {
    int32_t b;
  };
};

cell tSingle single {
};
