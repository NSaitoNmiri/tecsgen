/*
 * �ʲ����Զ���ƥ��Ȥ�����Ū�Ǻ��� 
 * Makefile �Ǥ� -U ����ꤹ��
 * 
 * [�Զ��] #516 ̾���ʤ� require �δؿ���¾�θƤӸ��δؿ�̾�Ƚ�ʣ�������ĸ�Ԥ���Ŭ������ʤ��ȡ�����ѥ�������顼
 * [�Զ��] #515 ��Ŭ���ʤ� -U �� require �ƤӸ��ν�ǥ���ѥ�������顼
 *                �ؿ�̾�� "__T" ����֤��뤳�Ȥǲ��
 */
signature sSig {
	int func( void );
};

/* Required Celltype & Cell */
[singleton]
celltype tRequired {
	entry sSig eEnt;
};
cell tRequired Required {
};

[singleton]
celltype tCelltype {
	require Required.eEnt;
	call    sSig     cCall;
};

cell tCelltype Cell {
	cCall = Required.eEnt;
};
