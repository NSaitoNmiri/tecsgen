/*
 * simple �ʥ���ץ�
 *
 * ���Υ���ץ�� tecsgen/test/simple ���ؤ��֤��Ƽ¹Ԥ���
 * Linux, Cygwin �Ķ��Ǽ¹ԤǤ���Ϥ�
 */

import_C( "tecs.h" );
import( <cygwin_kernel.cdl> );
import( <tSysLog.cdl> );

/* SysLog */
cell tSysLog SysLog {};

/* Kernel */
cell tKernel Kernel {};

/* typedef int32_t ER; */

signature sSimple {
	ER  func1( [in]int32_t inval );
	ER  func2( [out,string]char_t *str );
};

celltype tSimpleServer {
	entry sSimple eEnt;
};

celltype tSimpleClient {
	call sSimple cCall;
};

cell tSimpleServer SimpleServer {
};

cell tSimpleClient SimpleClient {
	[through(TracePlugin,"")]
		cCall = SimpleServer.eEnt;
};
