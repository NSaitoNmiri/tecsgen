/*
 *  TECS Generator
 *      Generator for TOPPERS Embedded Component System
 *  
 *   Copyright (C) 2008-2013 by TOPPERS Project
 *--
 *   �嵭����Ԥϡ��ʲ���(1)(4)�ξ������������˸¤ꡤ�ܥ��եȥ���
 *   �����ܥ��եȥ���������Ѥ�����Τ�ޤࡥ�ʲ�Ʊ���ˤ���ѡ�ʣ������
 *   �ѡ������ۡʰʲ������ѤȸƤ֡ˤ��뤳�Ȥ�̵���ǵ������롥
 *   (1) �ܥ��եȥ������򥽡��������ɤη������Ѥ�����ˤϡ��嵭������
 *       ��ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ��꤬�����Τޤޤη��ǥ���
 *       ����������˴ޤޤ�Ƥ��뤳�ȡ�
 *   (2) �ܥ��եȥ������򡤥饤�֥������ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ�����Ǻ����ۤ�����ˤϡ������ۤ�ȼ���ɥ�����ȡ�����
 *       �ԥޥ˥奢��ʤɡˤˡ��嵭�����ɽ�����������Ѿ�浪��Ӳ���
 *       ��̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *   (3) �ܥ��եȥ������򡤵�����Ȥ߹���ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ��ʤ����Ǻ����ۤ�����ˤϡ����Τ����줫�ξ�����������
 *       �ȡ�
 *     (a) �����ۤ�ȼ���ɥ�����ȡ����Ѽԥޥ˥奢��ʤɡˤˡ��嵭����
 *         �ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *     (b) �����ۤη��֤��̤�������ˡ�ˤ�äơ�TOPPERS�ץ������Ȥ�
 *         ��𤹤뤳�ȡ�
 *   (4) �ܥ��եȥ����������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������뤤���ʤ�»
 *       ������⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ����դ��뤳�ȡ�
 *       �ޤ����ܥ��եȥ������Υ桼���ޤ��ϥ���ɥ桼������Τ����ʤ���
 *       ͳ�˴�Ť����ᤫ��⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ�
 *       ���դ��뤳�ȡ�
 *  
 *   �ܥ��եȥ������ϡ�̵�ݾڤ��󶡤���Ƥ����ΤǤ��롥�嵭����Ԥ�
 *   ���TOPPERS�ץ������Ȥϡ��ܥ��եȥ������˴ؤ��ơ�����λ�����Ū
 *   ���Ф���Ŭ������ޤ�ơ������ʤ��ݾڤ�Ԥ�ʤ����ޤ����ܥ��եȥ���
 *   �������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������������ʤ�»���˴ؤ��Ƥ⡤��
 *   ����Ǥ�����ʤ���
 *  
 *   $Id: RPCTask.cdl 1925 2013-01-20 05:55:58Z okuma-top $
 */

/*
 * unmarshaler �� main �Υ����˥���
 */
signature sUnmarshalerMain {
	ER	main(void);
};

///////////////// ��ͭ�����ͥ��Ѥ���� ////////////////
/*
 * CELLTYPE: ��ͭ�����ͥ��ѤΥ������ᥤ��
 */
celltype tRPCDedicatedTaskMain {			// Transparent RPC ���Ѥ���
	entry	sTaskBody			eMain;
	call	sUnmarshalerMain	cMain;
};

celltype tRPCDedicatedTaskMainWithOpener {	// Opaque RPC ���Ѥ���
	entry	sTaskBody				eMain;
	call	sUnmarshalerMain		cMain;
	call	sServerChannelOpener	cOpener;
	attr {
		RELTIM	initialDelay = 0;	// sec
		RELTIM	reopenDelay = 1;	// sec
	};
	require tKernel.eKernel;
};

///////////////// ��ͭ�����ͥ��Ѥ���� ////////////////
/*
 * CONST: ��ͭ�����ͥ�إå��Υޥ��å�
 */
const uint16_t RPC_CHANNEL_MAN_SOP_MAGIC   = (0x3141);  // Beginning of using shared channel
const uint16_t RPC_CHANNEL_MAN_EOP_MAGIC   = (0x2718);  // End of using shared channel

/*
 * CELLTYPE: ��ͭ�����ͥ�ޥ͡�����
 * REM:      �ƤӸ�¦���֤������ͥ�ޥ͡�����
 *           eSemaphore ���ƤӽФ��줿�Ȥ������ͥ���å�����ȤȤ�ˡ�
 *           �����ͥ��ֹ�����Ф���
 */
celltype tRPCSharedChannelMan {
	entry	sSemaphore	eSemaphore[];
	call	sSemaphore	cSemaphore;
	call	sTDR		cClientSideTDR;
};


/*
 * CELLTYPE: ��ͭ�����ͥ��ѤΥ������ᥤ��
 * REM:      �Ƥ���¦���֤�������
 *           �����ͥ��ֹ����Ф��������ͥ��ֹ�� cTaskBody ��ƤӽФ�
 */
celltype tRPCSharedTaskMain {
	entry	sTaskBody	eMain;

	call	sUnmarshalerMain	cUnmarshalAndCallFunction[];
	call	sTDR		cServerSideTDR;

	require	tSysLog.eSysLog;

	var {
		int16_t	channelNo;	/* ����ź�� + 1 */
	};
};

celltype tRPCSharedTaskMainWithOpener {	// Opaque RPC ���Ѥ���
	entry	sTaskBody			eMain;
	call	sUnmarshalerMain	cUnmarshalAndCallFunction[];
	call	sTDR				cServerSideTDR;
	call	sServerChannelOpener cOpener;
	require	tSysLog.eSysLog;
	require tKernel.eKernel;

	attr {
		RELTIM	initialDelay = 0;	// sec
		RELTIM	reopenDelay = 1;	// sec
	};
	var {
		int16_t	channelNo;	/* ����ź�� + 1 */
	};
};
