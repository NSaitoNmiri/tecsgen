import_C( "tecs.h" );
import_C( "mydef.h" );
import( <cygwin_kernel.cdl> );
import( <tSysLog.cdl> );

cell tSysLog SysLog{};
cell tKernel Kernel{};

// typedef int32_t ER;

signature sSig1 {
	ER		func1( [in]int32_t a );
	int32_t	func2( [in]int32_t a );
};

signature sSig2 {
	ER		func1( [in]int32_t a );
	int32_t	func2( [in]int32_t a );
};

signature sSig3 {
	ER		func1( [in]int32_t a );
	int32_t	func2( [in]int32_t a );
};

celltype tCell1 {
	call sSig1 cCall;
	entry sSig2 eEntry;
	attr {
		int32_t a = C_EXP( "VAL_$id$" );
	};
	var {
		int32_t b = a;
	};
};

celltype tCell2 {
	call sSig2 cCall;
	entry sSig3 eEntry;
	attr {
		int32_t a;
		int32_t b = 10;
	};
	var {
		int32_t c[2] = { 1, 2 };
	};
};

composite tComposite {

	call	sSig1	cCall1;
	entry	sSig3	eEntry;
	attr {
		int32_t a = 100;
		int32_t b = C_EXP( "VAL_$id$" );
	};

	cell tCell1 cell1 {
		a = composite.a;
		cCall => composite.cCall1;
	};

	cell tCell2 cell2 {
		a = composite.a;
		b = composite.b;
		cCall = cell1.eEntry;
	};
	composite.eEntry => cell2.eEntry;
};

celltype tCell_serv{
	entry	sSig1	eEntry;
	attr {
		int32_t a;
	};
};

[singleton,active]
celltype tCell_clnt {
	call	sSig3	cCall;
	attr {
		int32_t a;
	};
};

cell tCell_serv cell_serv{
	a = 5;
};

cell tComposite compcell1 {
	// a=10;
	a = C_EXP( "VAL_$id$" );
	cCall1 = cell_serv.eEntry;
};

cell tComposite compcell2 {
	/* a=20; */
	cCall1 = cell_serv.eEntry;
};

cell tCell_clnt cell_clnt {
	a = 30;
	cCall = compcell1.eEntry;
};



[active,singleton]
celltype tCell2_active_single {
	call	sSig2	cCall;
	entry	sSig3	eEntry;
	attr {
		int32_t a;
	};
	var {
		int32_t b;
	};
};

[active,singleton]
composite tComposite_active_singleton {

	attr {
		int32_t	a = 2000;
	};
	call	sSig1	cCall1;
	entry	sSig3	eEntry;

	cell tCell1 cell1 {
		a = composite.a;
		cCall => composite.cCall1;
	};

	cell tCell2_active_single cell2 {
		a = composite.a;
		cCall = cell1.eEntry;
	};
	eEntry => cell2.eEntry;
};

cell tCell_serv cell_serv2{
	a = 5;
};
cell tComposite_active_singleton active_singleton {
	/* a = 30; */
	cCall1 = cell_serv2.eEntry;
};


int8_t * const PTRVAL = (int8_t *)0x1000;
//int8_t * const PTRVAL = 0x1000;

[active]
celltype tPtrAttr {
	attr {
		int8_t *p_attr0;
		int8_t *p_attr1;
		int8_t *p_attr2;
		int8_t *p_attr3 = (int8_t *)0x10;
	};
};

[active]
composite tCompPtrAttr {
	attr{
		int8_t *p_attr0;
		int8_t *p_attr1 = (int8_t *)0x20;
	};
	cell tPtrAttr PtrAttr{
		p_attr0 = composite.p_attr0;
		p_attr1 = composite.p_attr1;
		p_attr2 = (int8_t *)0x40;
	};
};

cell tCompPtrAttr PtrAttr {
	p_attr0 = (int8_t *)0x50;
};

cell tCompPtrAttr PtrAttr2 {
//	p_attr0 = (int8_t *)PTRVAL;
	p_attr0 = PTRVAL;
};

celltype tSizeArray {
	attr {
		int32_t  size;
		[size_is(size)]
			int8_t  *array;
	};
	factory {
		write( "tSizeArray.cfg", "tSizeArray: $id$" );
	};
};

cell tSizeArray SizeArray {
	size = 2;
	array = { 0, 1 };
};

composite tCompSizeArray {
	attr {
		int32_t siz;
		[size_is(siz)]
			int8_t *array;  // #386 �ǥ��顼�Ȥ���, #418 ����Ǥ褤����
	};
	cell tSizeArray Cell{
		size = composite.siz;
		array = composite.array;
	};
};

cell tCompSizeArray CompSizeArray {
	siz = 5;
	array = { 0 };    // #386 �㳰ȯ��
};


[active]
composite tOuterCompPtrAttr {
	attr{
		int8_t *p_attr0;
		int8_t *p_attr1;
	};
	cell tCompPtrAttr PtrAttr{
		p_attr0 = composite.p_attr0;
		p_attr1 = composite.p_attr1;
	};
};

/* �����ƤӸ��˹�ή���� */
composite tComp {
	call sSig1 cCall;
	cell tCell1 CellA {
		cCall => composite.cCall;
	};
	cell tCell1 CellB {
		cCall => composite.cCall;
	};
};

//	[through(TracePlugin,"")]
