/*
 * simple �ʥ���ץ�
 *
 * ���Υ���ץ�� tecsgen/test/simple ���ؤ��֤��Ƽ¹Ԥ���
 * Linux, Cygwin �Ķ��Ǽ¹ԤǤ���Ϥ�
 *
 * tecs_package for OpaqueRPC �Ȱ��פ����Ƥ���
 */
import_C( "cygwin_tecs.h" );
import_C( "my_setjmp.h" );

// ����ǽ
import( <tSysLog.cdl> );
// �����ͥ뵡ǽ
import( <cygwin_kernel.cdl> );
import( <rpc.cdl> );
import( <tSocketChannel.cdl> );
import( "tAlloc.cdl" );
import( "sSimple.cdl" );

/// Server Celltype ///
celltype tSimpleServer {
	require	tSysLog.eSysLog;
	entry	sSimple			eEnt;
/*	entry	sServerControl	eServerControl; */
};

/// Client Celltype ///
[active]
celltype tSimpleClient {
	require	tSysLog.eSysLog;
	call	sSimple		cCall;
	/* call	sServerControl	cServerControl;	/* �����Ф򥷥�åȥ����󤹤� */
	call	sSocketClientOpener	cOpener;	/* �����ͥ�򳫤� */
	entry	sTaskBody	eMain;					/* �ᥤ�� */
	entry   sRPCErrorHandler eHandler;
	var {
		jmp_buf  jbuf;
	};
};

/// Error Handler Celltype Client side & Server side ///
celltype tClientRPCErrorHandler {
	entry sRPCErrorHandler eHandler;
	call sRPCErrorHandler cHandler;
};
celltype tServerRPCErrorHandler {
	entry sRPCErrorHandler eHandler;
	call  sServerChannelOpener cOpener;
};

// to_through �ǻ��ѤǤ��뤽��¾�Υ��ץ���� ( '\"', '%', '!' ���Ȥ��� )��
//			"clientChannelCelltype= "\tSocketClient"\, "		// ���饤�����¦�����ͥ륻�륿����̾
//			"serverChannelCelltype= "\tSocketClient"\, "		// �����С�¦�����ͥ륻�륿����̾
//			"clientChannelInitializer= !portNo=8931+$count$; serverAddr=\"127.0.0.1\";!, "
//			"serverChannelInitializer= !portNo=8931+$count$;!, "	// �����ͥ�
//			"clientSemaphoreInitializer= !count = 1; attribute = C_EXP( \"TA_NULL\" );! ,"
//			"clientSemaphoreCelltype = tCelltype;, "                // ���ޥե����륿����
//			"TDRCelltype=\"tNBOTDR\","
//			"taskCelltype=tTask,"									// �����С�¦���������륿����
//			"taskPriority=11,"										// �����С�¦������ͥ����
//			"StackSize=4096,"										// �����С�¦�����������å�������
//  ���Ū�Τ��ᡢ'!', '%', "'", "\"" ��ȤäƤ��뤬���ɤ�Ǥ�Ʊ���Ǥ��롣
//  ����������������� \" ��Ȥ��������ˤϡ�����ʳ�����Ѥ���ɬ�פ����롣
//  �֤� ',' ���ʤ��ΤǤ���С�ɬ�����⡢�����ǳ��ɬ�פϤʤ���

//[ out_through(),   out_through �����פˤʤä�  V1.B.0.11
[to_through(rServer ,OpaqueRPCPlugin,
			"PPAllocatorSize=1024,"									// PPAllocator ������(����������)
			"substituteAllocator=%Alloc.eAlloc=>CAlloc.eAlloc%, "	// ���إ����������� (�ǥե���Ȥ�̤����)
			"clientChannelCell= 'ClientChannel_$destination$', "	// ���饤�����¦�����ͥ륻��̾
			"serverChannelCell= !ServerChannel_$destination$!,  "	// �����С�¦�����ͥ륻��̾
			"clientErrorHandler = 'ClientRPCErrorHandler_$destination$.eHandler', " // ���顼�ϥ�ɥ顼 (�ǥե���Ȥ�̤����)
			"serverErrorHandler = 'ServerRPCErrorHandler_$destination$.eHandler', " // ���顼�ϥ�ɥ顼 (�ǥե���Ȥ�̤����)
//			"clientChannelInitializer= !portNo=8931+$count$; serverAddr=\"192.168.99.1\";!, "
				//  cygwin �Υ��饤����Ȥ� skyeye �Υ����С�����³���ƻ����ݤ�����
				//  README-skyeyeWithTINET.pdf �򻲾ȤΤ���
			), linkunit]
region rClient /*,nNamespace */ {
	cell tSysLog ClientSysLog {
	};
	cell tAlloc CAlloc {
	};
	cell tKernel KernelInClient {
	};

	// RPC Error Handler Client Side
	cell tClientRPCErrorHandler ClientRPCErrorHandler_SimpleServer{
		cHandler = rCPon::SimpleClient.eHandler;
	};

	// [out_through(TracePlugin,""),in_through()]
	[out_through(),in_through()]
	region rCPon {
		cell tSimpleClient SimpleClient {
			[through(TracePlugin,"")]
				cCall = rServer::rSPon::SimpleServer.eEnt;
			cOpener = ClientChannel_SimpleServer.eOpener;
		};
		cell tTask Task {
			cBody = SimpleClient.eMain;
			priority = 1;
			stackSize = 4096;
			taskAttribute = C_EXP( "TA_ACT" );
		};
	};
};

[linkunit]
region rServer {
	cell	tSysLog	ServerSysLog {
	};
	cell tKernel KernelInServer {
	};
	// RPC Error Handler Server Side
	cell tServerRPCErrorHandler ServerRPCErrorHandler_SimpleServer{
		cOpener = ServerChannel_SimpleServer.eOpener;
	};

	[in_through(TracePlugin,""),out_through()]
		// [in_through()]
	region rSPon {
    //      cell tSysLog ServerSysLog {
    //      };
		cell tAlloc Alloc {
		};
		[allocator(eEnt.func21.a=Alloc.eAlloc,
				   eEnt.func22.sta=Alloc.eAlloc,
				   eEnt.func23.str=Alloc.eAlloc,
				   eEnt.func24.msg=Alloc.eAlloc,
				   eEnt.func25.msg=Alloc.eAlloc,
				   eEnt.func26.sta=Alloc.eAlloc,
				   eEnt.func27.array2=Alloc.eAlloc,
				   eEnt.func31.a=Alloc.eAlloc,
				   eEnt.func32.sta=Alloc.eAlloc,
				   eEnt.func33.str=Alloc.eAlloc,
				   eEnt.func34.msg=Alloc.eAlloc,
				   eEnt.func35.msg=Alloc.eAlloc,
				   eEnt.func36.sta=Alloc.eAlloc,
				   eEnt.func37.sta=Alloc.eAlloc,
				   eEnt.func38.array2=Alloc.eAlloc,
				   eEnt.func39.arraySt=Alloc.eAlloc)]
		cell tSimpleServer SimpleServer {
		};
	};
};

