/*
 * ��require�ƥ��ȥ�����
 *
 * �ʲ���4�ĤΥ�������ƥ��Ȥ���
 * (1) ���륿���פ� entry �ǵ�require (celltype) �����ꤵ��Ƥ��� (ɸ��Ū�ʻȤ���)
 * (2) ���륿���פ� entry �ǵ�require (cell) �����ꤵ��Ƥ��� (ɸ��Ū�ʻȤ���)
 * (3) composite �������Υ���˵�require�����ꤵ��Ƥ���
 * (4) composite �� entry �ǵ�require�����ꤵ��Ƥ���
 *
 * �����Υƥ��ȥ������ˤϡ���require ���������̤η�礬�ʤ���Ƥ����2�İʾ�η�礬���뤳�ȡˤˤ�� warning ���Ф뤳�Ȥλ��Ԥ�
 */

import_C( "cygwin_tecs.h" );

signature sInit {
	void initialize( void );
};

[singleton,active]
celltype tInitializer {
   call sInit cInit[];
};

cell tInitializer Initializer {
	cInit[] = Cell11.eInit;      /* �� require ���ꤵ��Ƥ��륻�� (warning) */
	cInit[] = Cell21.eInit;      /* �� require ���ꤵ��Ƥ��륻�� (warning) */
	cInit[] = CompCell31.eInit;  /* �� require ���ꤵ��Ƥ��륻�� (warning) */
	cInit[] = CompCell41.eInit;  /* �� require ���ꤵ��Ƥ��륻�� (warning) */
	cInit[] = CompCell51.eInit;  /* �� require ���ꤵ��Ƥ��륻�� (warning) */
};

// (1) ��require �򥻥륿���פǻ��ꤹ����
celltype tCelltype {
	// entry sInit eInit <= Initializer.cInit;
	entry sInit eInit <= tInitializer.cInit;
	attr {
		int32_t  no;
	};
};

cell tCelltype Cell11 {
	no = 11;
};


cell tCelltype Cell12 {
	no = 12;
};


// (2) ��require �򥻥�ǻ��ꤹ����
celltype tCelltype2 {
	entry sInit eInit <= Initializer.cInit;
	// entry sInit eInit <= tInitializer.cInit;
	attr {
		int32_t  no;
	};	
};


cell tCelltype2 Cell21 {
	no = 21;
};


cell tCelltype2 Cell22 {
	no = 22;
};

/* (3) composite ���륿���פ���¦�Υ���ǡ��� require �����ꤵ��Ƥ��� */
composite tComposite {
	attr{ int32_t no; };
	entry sInit eInit;       /* ��requie ���ꤵ��Ƥ���������� export */
	cell tCelltype2 Cell {
		no = composite.no;
	};
	composite.eInit => Cell.eInit;
};

cell tComposite CompCell31 {
	no = 31;
};

cell tComposite CompCell32 {
	no = 32;
};

// (4) ��require �򥻥�ǻ��ꤹ����
celltype tCelltype3 {
	entry sInit eInit;
	attr {
		int32_t  no;
	};	
};

/* (4-1) composite ���륿���פ� entry �ǡ��� require �����ꤵ��Ƥ��� */
composite tComposite2 {
	entry sInit eInit <= tInitializer.cInit;
	attr {
		int32_t no;
	};

	cell tCelltype3 Cell {
		no = composite.no;
	};
	composite.eInit => Cell.eInit;
};

/* (4-2) */
composite tComposite3 {
	entry sInit eInit <= Initializer.cInit;
	attr {
		int32_t no;
	};

	cell tCelltype3 Cell {
		no = composite.no;
	};
	composite.eInit => Cell.eInit;
};

cell tComposite2 CompCell41 {
	no = 41;
};

cell tComposite3 CompCell42 {
	no = 42;
};

composite tCompositeOuter {
	entry sInit eInit;
	attr {
		int32_t no;
	};

	cell tComposite Cell {
		no = composite.no;
	};
	composite.eInit => Cell.eInit;
};

cell tCompositeOuter CompCell51 {
	no = 51;
};
