typedef int32_t ER;

signature sSyscall{
	ER func( void );
};

signature sSyscall2{
	ER func( void );
};

[singleton]
celltype tKernel {
	entry sSyscall eSc;
	entry sSyscall2 eSc2;
};
cell tKernel Kernel {
};

/* require �ǥ���̾����� */
celltype tRequire{
	require Kernel.eSc;
	require Kernel.eSc2;
};

cell tRequire Require {
};


/* require �ǥ��륿����̾����� */
celltype tRequire2{
	require tKernel.eSc;
	require tKernel.eSc;
};

cell tRequire2 Require2 {
};
