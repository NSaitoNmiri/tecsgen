/* �꡼����󤴤Ȥ˥����ɤ���������ƥ��� */
/* tecsgen -G rRegion2 �ˤ�� rRegion2 �Τ߽��� */

import_C( "tecs.h" );

/* typedef int32_t ER; */

signature sMain {
	void  main(void);
};

signature sSig1 {
	ER func1( [in]int32_t arg1, [out]int32_t *res );
};

signature sSig2 {
	ER func1( [in]int32_t arg1, [out]int32_t *res );
};

signature sSig3 {
	ER func1( [in]int32_t arg1, [out]int32_t *res );
};

celltype tCtR1 {
	entry sSig3 eEnt;
};

celltype tCtR2 {
	call sSig2 cCall2;
	call sSig3 cCall3;
	entry sSig1 eEnt;
};

celltype tCtOuter {
	call    sSig1  cCall;
	entry   sSig2  eEnt;
	entry   sMain  eMain;
	attr{
		int32_t  a;
	};
};

[singleton]
celltype tSingle {
	attr {
		int32_t  Attr;
	};
};

/* rRegion2 ��и��� specifier ����� */
[to_through(rRegion1, TracePlugin, ""),
out_through(/*TracePlugin,""*/),
in_through()]
region rRegion2 {
	/* �ץ�ȥ�������� */
	cell tCtR2 r2cell;
};

/* rRegion1 ��и��� specifier ����� */
[in_through(/*TracePlugin, ""*/)]
region rRegion1{
	/* �ץ�ȥ�������� */
	cell tCtR1 r1cell;
};

cell tCtOuter outer {
	cCall = rRegion2::r2cell.eEnt;
	a = 0;
};

/* �����ʺƽи��ˤǤ� specifier �����Ǥ��ʤ� */
region rRegion1 {
	cell tCtR1 r1cell {
	};
	cell tSingle Single1 {
		Attr = 10;
	};
};

/* �����ʺƽи��ˤǤ� specifier �����Ǥ��ʤ� */
region rRegion2 {
	cell tCtOuter outer2 {
		cCall = r2cell.eEnt;
		a = 101;
	};

	cell tCtR1 r1cell2 {
	};
	cell tCtR2 r2cell {
		cCall2 = outer2.eEnt;
		cCall3 = r1cell2.eEnt;
	};

	[out_through()]
	region rRegionInner {
		cell tCtR2 r2cellInner {
			cCall2 = outer.eEnt;
			cCall3 = r1cell2.eEnt;
		};
	};
};

[singleton,active]
celltype tMain {
	call sMain cMain;
};

region rRegion2 {
	cell tMain Main{
		cMain = outer2.eMain;
	};

	/* 2���ܤ� tSingle */
//	cell tSingle Single2 {
//		Attr = -999;
//	};
};

