const int32_t consVal = C_EXP( "AA" );
const int32_t consVal2 = consVal;

celltype tC_exp {
	attr {
		int32_t id = C_EXP( "ID_$id$" );
		char_t *cbp = C_EXP( "\"cell: $cell$, ct: $ct$, idx: $idx$, cb_proto: $cb_proto$, cbp: $cbp$, id: $id$\"\n" );
	};
	var {
		int32_t v = C_EXP( "false" );
	};
	factory{
		write( "tecsgen.cfg", "CRE_SEM(SEMID_SERIALPORT_$id$_SND,  { TA_TPRI, 0, 1 })" );
		write( "tecsgen.cfg", "cbp:: \"%s\"", cbp );
		write( "tecsgen.cfg", "cbp:: %s", cbp );
		write( "tecsgen.cfg", "id:: %s\n", id );
	};
};

cell tC_exp tc {
};

// composite $B$N>l9g(B
// $cell$, $id$, $ct$ $B$O!"(Bcomposite $B%;%k$N$b$N$H$J$k!JFbIt%;%k$N$b$N$O;H$o$l$J$$!K(B
// $idx$, $cb_proto$, $cbp$ $B$O<BBN$KBP$9$k$b$N$J$N$G!"FbIt%;%k$N$b$N$H$J$k(B
composite tComp_C_EXP {
	attr {
		char_t *cbp = C_EXP( "\"cell: $cell$, ct: $ct$, idx: $idx$, cb_proto: $cb_proto$, cbp: $cbp$, id: $id$\"" );
	};
	cell tC_exp tc {
		cbp = composite .cbp;
		id = C_EXP( "\"ID_$id$_CELL_$cell$_IDX_$idx$, CB_PROTO $cb_poroto$, CBP $cbp$\"" );
	};
};

cell tComp_C_EXP tc2 {
};

cell tComp_C_EXP tc3 {
	cbp =  C_EXP( "\"TC3: cell: $cell$, ct: $ct$, idx: $idx$, cb_proto: $cb_proto$, cbp: $cbp$, id: $id$\"" );
};
