/*
 *  TECS Generator
 *      Generator for TOPPERS Embedded Component System
 *  
 *   Copyright (C) 2008-2013 by TOPPERS Project
 *--
 *   �嵭����Ԥϡ��ʲ���(1)(4)�ξ������������˸¤ꡤ�ܥ��եȥ���
 *   �����ܥ��եȥ���������Ѥ�����Τ�ޤࡥ�ʲ�Ʊ���ˤ���ѡ�ʣ������
 *   �ѡ������ۡʰʲ������ѤȸƤ֡ˤ��뤳�Ȥ�̵���ǵ������롥
 *   (1) �ܥ��եȥ������򥽡��������ɤη������Ѥ�����ˤϡ��嵭������
 *       ��ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ��꤬�����Τޤޤη��ǥ���
 *       ����������˴ޤޤ�Ƥ��뤳�ȡ�
 *   (2) �ܥ��եȥ������򡤥饤�֥������ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ�����Ǻ����ۤ�����ˤϡ������ۤ�ȼ���ɥ�����ȡ�����
 *       �ԥޥ˥奢��ʤɡˤˡ��嵭�����ɽ�����������Ѿ�浪��Ӳ���
 *       ��̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *   (3) �ܥ��եȥ������򡤵�����Ȥ߹���ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ��ʤ����Ǻ����ۤ�����ˤϡ����Τ����줫�ξ�����������
 *       �ȡ�
 *     (a) �����ۤ�ȼ���ɥ�����ȡ����Ѽԥޥ˥奢��ʤɡˤˡ��嵭����
 *         �ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *     (b) �����ۤη��֤��̤�������ˡ�ˤ�äơ�TOPPERS�ץ������Ȥ�
 *         ��𤹤뤳�ȡ�
 *   (4) �ܥ��եȥ����������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������뤤���ʤ�»
 *       ������⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ����դ��뤳�ȡ�
 *       �ޤ����ܥ��եȥ������Υ桼���ޤ��ϥ���ɥ桼������Τ����ʤ���
 *       ͳ�˴�Ť����ᤫ��⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ�
 *       ���դ��뤳�ȡ�
 *  
 *   �ܥ��եȥ������ϡ�̵�ݾڤ��󶡤���Ƥ����ΤǤ��롥�嵭����Ԥ�
 *   ���TOPPERS�ץ������Ȥϡ��ܥ��եȥ������˴ؤ��ơ�����λ�����Ū
 *   ���Ф���Ŭ������ޤ�ơ������ʤ��ݾڤ�Ԥ�ʤ����ޤ����ܥ��եȥ���
 *   �������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������������ʤ�»���˴ؤ��Ƥ⡤��
 *   ����Ǥ�����ʤ���
 *  
 *   $Id: $
 */


/* client side state */
const	int16_t	RPCSTATE_CLIENT_GET_SEM		= 1;
const	int16_t	RPCSTATE_CLIENT_SEND_SOP	= 2;
const	int16_t	RPCSTATE_CLIENT_SEND_BODY	= 3;
const	int16_t	RPCSTATE_CLIENT_SEND_EOP	= 4;
const	int16_t	RPCSTATE_CLIENT_EXEC		= 5;
const	int16_t	RPCSTATE_CLIENT_RECV_SOP	= 6;
const	int16_t	RPCSTATE_CLIENT_RECV_BODY	= 7;
const	int16_t	RPCSTATE_CLIENT_RECV_EOP	= 8;
const	int16_t	RPCSTATE_CLIENT_RELEASE_SEM	= 9;

/* server side state */
const	int16_t	RPCSTATE_SERVER_GET_SEM		= 11;
const	int16_t	RPCSTATE_SERVER_RECV_SOP	= 12;
const	int16_t	RPCSTATE_SERVER_RECV_BODY	= 13;
const	int16_t	RPCSTATE_SERVER_RECV_EOP	= 14;
const	int16_t	RPCSTATE_SERVER_EXEC		= 15;
const	int16_t	RPCSTATE_SERVER_SEND_SOP	= 16;
const	int16_t	RPCSTATE_SERVER_SEND_BODY	= 17;
const	int16_t	RPCSTATE_SERVER_SEND_EOP	= 18;
const	int16_t	RPCSTATE_SERVER_RELEASE_SEM	= 19;

/* error hadler */
signature sRPCErrorHandler {
	ER	errorOccured( [in]int16_t func_id, [in]ER er, [in]int16_t state );
};

/*
 * �ƤӸ�¦�Ǥ� state �� RPCSTATE_CLIENT_EXEC �����������礭����硢
 * �Ƥ���¦�Ǥ� state �� RPCSTATE_SERVER_EXEC �����������礭����硢
 * �Ƥ���ؿ��θƤӽФ��ˤ��������Ƥ��롣
 *
 * RPCErrorHandler ���ƤӽФ��줿�����ǡ�send/receive �����β����Ͻ���äƤ��롣
 * ���Τ��ᡢRPCErrorHandler ����ǽ������Ǥ��ڤäƤ�(�������κƵ�ư�ʤɤ�ԤäƤ�)�������ˤ�����꡼���������ʤ���
 */
