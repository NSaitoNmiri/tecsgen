/*
 *  TECS Generator
 *      Generator for TOPPERS Embedded Component System
 *  
 *   Copyright (C) 2008-2013 by TOPPERS Project
 *--
 *   �嵭����Ԥϡ��ʲ���(1)(4)�ξ������������˸¤ꡤ�ܥ��եȥ���
 *   �����ܥ��եȥ���������Ѥ�����Τ�ޤࡥ�ʲ�Ʊ���ˤ���ѡ�ʣ������
 *   �ѡ������ۡʰʲ������ѤȸƤ֡ˤ��뤳�Ȥ�̵���ǵ������롥
 *   (1) �ܥ��եȥ������򥽡��������ɤη������Ѥ�����ˤϡ��嵭������
 *       ��ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ��꤬�����Τޤޤη��ǥ���
 *       ����������˴ޤޤ�Ƥ��뤳�ȡ�
 *   (2) �ܥ��եȥ������򡤥饤�֥������ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ�����Ǻ����ۤ�����ˤϡ������ۤ�ȼ���ɥ�����ȡ�����
 *       �ԥޥ˥奢��ʤɡˤˡ��嵭�����ɽ�����������Ѿ�浪��Ӳ���
 *       ��̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *   (3) �ܥ��եȥ������򡤵�����Ȥ߹���ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ��ʤ����Ǻ����ۤ�����ˤϡ����Τ����줫�ξ�����������
 *       �ȡ�
 *     (a) �����ۤ�ȼ���ɥ�����ȡ����Ѽԥޥ˥奢��ʤɡˤˡ��嵭����
 *         �ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *     (b) �����ۤη��֤��̤�������ˡ�ˤ�äơ�TOPPERS�ץ������Ȥ�
 *         ��𤹤뤳�ȡ�
 *   (4) �ܥ��եȥ����������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������뤤���ʤ�»
 *       ������⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ����դ��뤳�ȡ�
 *       �ޤ����ܥ��եȥ������Υ桼���ޤ��ϥ���ɥ桼������Τ����ʤ���
 *       ͳ�˴�Ť����ᤫ��⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ�
 *       ���դ��뤳�ȡ�
 *  
 *   �ܥ��եȥ������ϡ�̵�ݾڤ��󶡤���Ƥ����ΤǤ��롥�嵭����Ԥ�
 *   ���TOPPERS�ץ������Ȥϡ��ܥ��եȥ������˴ؤ��ơ�����λ�����Ū
 *   ���Ф���Ŭ������ޤ�ơ������ʤ��ݾڤ�Ԥ�ʤ����ޤ����ܥ��եȥ���
 *   �������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������������ʤ�»���˴ؤ��Ƥ⡤��
 *   ����Ǥ�����ʤ���
 *  
 *   $Id: PPAllocator.cdl 1925 2013-01-20 05:55:58Z okuma-top $
 */

/*
 * PPAlloc: Push Pop Allocator
 *
 * allocate �����ս�� deallocate ���ʤ��ƤϤʤ�ʤ�
 * deallocate �ϡ��ޤȤ�ƹԤ����Ȥ��Ǥ���
 * �㤨�кǽ�� allocate ���줿�ΰ�� deallocate ����ȡ����٤Ƥ� allocate ���줿�ΰ�� deallocate �������Ȥˤʤ�
 * ��¾���椷�Ƥ��ʤ�����ñ��Υ������˳��դ��ƻ��Ѥ���
 */

[deviate]   // alloc ����æ�ˤʤ�
signature sPPAllocator {
	/*
	 * size �ǻ��ꤵ�줿�礭���Υ����ΰ�򥢥����Ȥ���
	 * �����ΰ褬���ݤ��줿��� *ptr �˥����ΰ�Υ��ɥ쥹���Ǽ���� E_OK ���֤�
	 * ��ʬ�ʶ����ΰ褬�ʤ���� E_NOMEM ���֤�
	 */
	ER  alloc( [in]uint32_t size, [out]void **ptr );
	/*
	 * �����ǥ������Ȥ���
	 * alloc �ǳ��������ݥ��󥿤������ ptr �˻��ꤹ��
	 * alloc �ǳ������������ΰ�� alloc �����ΤȤϵս�� dealloc ���ʤ��ƤϤʤ�ʤ�
	 * ���٤Ƥ� dealloc ����ˤϡ��ǽ�� alloc ���줿�����ΰ�� dealloc ���뤳�ȤǹԤ����Ȥ��Ǥ���
	 * alloc ���������������ΰ�򤹤٤� dealloc �������ˡ��Ƥ� alloc ���뤳�ȤϤǤ���
	 * ���ξ��Ǥ⡢dealloc ���Ƥ��ʤ������ΰ�� alloc �����ΤȤϵս�� dealloc ���ʤ��ƤϤʤ�ʤ�
	 *
	 * ptr ���ͤ� buf <= ptr < buf+allocated_size �����������ɤ������������
	 * ptr ���ͤ������ξ�� E_PAR ���֤�
	 */
	ER  dealloc( [in]const void *ptr );

    /*
	 * PPAllocator ����γ��դ��Ѥߥ���򤹤٤Ʋ�������
	 * ���δؿ���ɬ����������
	 */
    ER  dealloc_all(void);
};

celltype tPPAllocator {
	entry  sPPAllocator ePPAllocator;
	attr {
		uint32_t   heapSize;
	};
	var {
		[size_is(heapSize)]
			int8_t  *buf;
		uint32_t   allocatedSize;
	};
};

