const float32_t   f_val = 1.0;              // ����
const float32_t   f_val2 = 1.0 << 2;        // ��ư������ << �Ǥ��ʤ�
const float32_t   f_val3 = 1 << 2.0;        // 2.0 ������ cast ��ɬ��
const double64_t  f_val4 = "abc";          // 
int16_t * const p = (int16_t *)"string";  // TECS �ǤϷ��Ѵ�������ʤ�
int16_t * const p = (int16_t *)1 << 32;   // pointer �ͤ򥷥եȤǤ��ʤ�
const int16_t  *p = (int16_t *)0xfff00;   // const �ǤϤʤ�
const int16_t   i_val1 = (int16_t)9999999999.999;   // �礭������
const int16_t   i_val2 = (int16_t)-9999999999.999;   // ����������
const uint16_t  i_val3 = (uint16_t)-9999999999.999;  // �����
const uint16_t  i_val4 = (uint16_t)-9999999999;      // ���������
const uint16_t  i_val5 = (uint16_t)-0xff123456;      // ���������
const uint16_t  i_val6 = "abc";          // 
const char_t  *const  p_str  = "abc";    // ����
const int8_t  *const  p_str1  = "abc";
const int16_t *const  p_str2  = "abc";
