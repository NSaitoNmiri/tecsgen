import( <posix.cdl> );

/*
 * tools/mruby/mruby.c $B$+$i(B cInit_initializeBridge( mrb ) $B$r8F$S=P$9$h$&$KJQ99$7$?$b$N(B
 */
namespace nMruby{
	[active]
	celltype tMrubyProc {
	    entry nPosix::sMain eMain;

		[optional]
			call sInitializeBridge cInit;
		var {
			mrb_state *mrb;
		};
	};
};
