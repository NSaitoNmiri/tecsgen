import_C( "cygwin_tecs.h" );
import("tSysLog.cdl" );
import("cygwin_kernel.cdl" );

/*
 * import �����ʤ����� plugin ��Ƥ�Ǥ�褤���Υƥ���
 * nest ���������ͥ졼���� region �� through ����äƽ��Ϥ��줿�ꡢ����ʤ��ä����ƥ���
 */

import( "region-body.cdl" );
