
celltype tAttribute6 {
	attr {
		int		*a = { 0, 1 };
	};
	var {
		int	*c = a;          /* $B=i4|CM$,(B { ... } */
	};
};

celltype tAttribute5 {
	attr {
		//		int		a = { 0, 1 };
		int		a = C_EXP( "a" );
		int		b = "abc";
	};
	var {
		[size_is(a)]          /* size_is $B$N0z?t$,(B C_EXP */
			int	*c;
		[size_is(b)]          /* size_is $B$N0z?t$,(B $BJ8;zNs(B */
			int	*d = a * 2;   /* C_EXP $B$NCM$r(B2$BG\$7$h$&$H$7$F$$$k(B */
	};
};

cell tAttribute5 Attribute5_1 {
	a = 2;
	b = 3;
};

cell tAttribute5 Attribute5_2 {
};
