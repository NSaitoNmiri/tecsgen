signature sSig {
  int32_t   func( void );
};

celltype tClient {
  call sSig cCall;
};
celltype tServer {
  entry sSig eEnt;
};

// [in_through()]
region rServer{
  cell tServer Server {
  };
};

/* in_through $B$G$-$J$$%1!<%9(B */
cell tClient Client {
	cCall = rServer::Server.eEnt;
};

// [out_through(), to_through(rNoOut,TracePlugin,"")]
// [out_through()]
region rClient{
  /* to_through $B$G$-$J$$%1!<%9(B */
  cell tClient Client {
     cCall = rServer::Server.eEnt;
  };
  /* out_through $B$G$-$J$$%1!<%9(B */
  cell tClient Client2 {
     cCall = Server.eEnt;
  };
};

cell tServer Server {
};
