/*
 *  TECS Generator
 *      Generator for TOPPERS Embedded Component System
 *  
 *   Copyright (C) 2008-2013 by TOPPERS Project
 *--
 *   �嵭����Ԥϡ��ʲ���(1)(4)�ξ������������˸¤ꡤ�ܥ��եȥ���
 *   �����ܥ��եȥ���������Ѥ�����Τ�ޤࡥ�ʲ�Ʊ���ˤ���ѡ�ʣ������
 *   �ѡ������ۡʰʲ������ѤȸƤ֡ˤ��뤳�Ȥ�̵���ǵ������롥
 *   (1) �ܥ��եȥ������򥽡��������ɤη������Ѥ�����ˤϡ��嵭������
 *       ��ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ��꤬�����Τޤޤη��ǥ���
 *       ����������˴ޤޤ�Ƥ��뤳�ȡ�
 *   (2) �ܥ��եȥ������򡤥饤�֥������ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ�����Ǻ����ۤ�����ˤϡ������ۤ�ȼ���ɥ�����ȡ�����
 *       �ԥޥ˥奢��ʤɡˤˡ��嵭�����ɽ�����������Ѿ�浪��Ӳ���
 *       ��̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *   (3) �ܥ��եȥ������򡤵�����Ȥ߹���ʤɡ�¾�Υ��եȥ�������ȯ�˻�
 *       �ѤǤ��ʤ����Ǻ����ۤ�����ˤϡ����Τ����줫�ξ�����������
 *       �ȡ�
 *     (a) �����ۤ�ȼ���ɥ�����ȡ����Ѽԥޥ˥奢��ʤɡˤˡ��嵭����
 *         �ɽ�����������Ѿ�浪��Ӳ�����̵�ݾڵ����Ǻܤ��뤳�ȡ�
 *     (b) �����ۤη��֤��̤�������ˡ�ˤ�äơ�TOPPERS�ץ������Ȥ�
 *         ��𤹤뤳�ȡ�
 *   (4) �ܥ��եȥ����������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������뤤���ʤ�»
 *       ������⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ����դ��뤳�ȡ�
 *       �ޤ����ܥ��եȥ������Υ桼���ޤ��ϥ���ɥ桼������Τ����ʤ���
 *       ͳ�˴�Ť����ᤫ��⡤�嵭����Ԥ����TOPPERS�ץ������Ȥ�
 *       ���դ��뤳�ȡ�
 *  
 *   �ܥ��եȥ������ϡ�̵�ݾڤ��󶡤���Ƥ����ΤǤ��롥�嵭����Ԥ�
 *   ���TOPPERS�ץ������Ȥϡ��ܥ��եȥ������˴ؤ��ơ�����λ�����Ū
 *   ���Ф���Ŭ������ޤ�ơ������ʤ��ݾڤ�Ԥ�ʤ����ޤ����ܥ��եȥ���
 *   �������Ѥˤ��ľ��Ū�ޤ��ϴ���Ū�������������ʤ�»���˴ؤ��Ƥ⡤��
 *   ����Ǥ�����ʤ���
 *  
 *   $Id: $
 */

import_C( "tecs_rpc.h" );

// Straight Order TDR
const uint32_t TDR_SOP_MAGIC1   = (0x672A);  // Client to Server
const uint32_t TDR_SOP_MAGIC2   = (0x561E);  // Server to Client
const uint32_t TDR_EOP_MAGIC1   = (0x5A3C);  // �ֿ����Ԥ� (Ʊ���ƽФ�)
const uint32_t TDR_EOP_MAGIC2   = (0x6D5E);  // �ֿ����Ԥ��ʤ�(��Ʊ���ƽФ��ޤ��ϥ꥿����)

// Straight Order TDR for SharedChannel
const uint32_t TDR_SHSOP_MAGIC1   = (0x98D5);  // Client to Server
const uint32_t TDR_SHSOP_MAGIC2   = (0xA9E1);  // Server to Client
const uint32_t TDR_SHEOP_MAGIC1   = (0xB5C3);  // �ֿ����Ԥ� (Ʊ���ƽФ�)
const uint32_t TDR_SHEOP_MAGIC2   = (0x92A1);  // �ֿ����Ԥ��ʤ�(��Ʊ���ƽФ��ޤ��ϥ꥿����)

/*
 * TDR: TECS Data Representation layer
 */
[deviate]         /* get_intptr ����æ�ˤʤ� */
signature sTDR {  /* TECS Data Representation */

	/* ����ؿ� */

	/* �����ͥ�Υꥻ�å� */
	ER	reset( void );	/* �̿������ͥ�Υꥻ�å� */
						/* ����ǥ��顼��ȯ�����������ޤ��ϼ�����³�ԤǤ��ʤ��ä��Ȥ��ϥꥻ�åȤ��� */
						/* �������ꥻ�åȤ򤫤���ȡ�¾���� RESET ���顼���֤� */
						/* ��ǧ�Ǥ��ʤ��Ȥ��ϡ����Υ���ͥ���������뤷���ʤ� */

	/* �ޥ��å������ɤ������� */
	ER	sendSOP( [in]bool_t b_client );     /* StartOfPacket magic ������ */
	ER	receiveSOP( [in]bool_t b_client );  /* StartOfPacket magic ����� */
						 /* b_client: ���饤�����¦�ʤ� true, �����С�¦�ʤ� false */

	/* �ޥ��å������ɤ������� */
	//	ER	sendSHSOP( [in]bool_t b_client );     /* StartOfPacket magic ������ */
	//	ER	receiveSHSOP( [in]bool_t b_client );  /* StartOfPacket magic ����� */
						 /* b_client: ���饤�����¦�ʤ� true, �����С�¦�ʤ� false */

	ER	sendEOP( [in]bool_t b_continue );   /* EndOfPacket magic �������ʥѥ��åȤ��ݤ�������Ԥ��� */
	ER	receiveEOP( [in]bool_t b_continue );/* EndOfPacket magic ����� */
                        /* b_continue: Ʊ���ƤӽФ��Υ��饤�����¦�ʤ� true,
                           ��Ʊ���ƤӽФ��Υ��饤�����¦�ޤ��ϥ����С�¦�ʤ� false */

	/* �ǡ����������ؿ� */

	/* ������ (�侩) */
	ER	putInt8( [in]int8_t in ); 
	ER	putInt16( [in]int16_t in ); 
	ER	putInt32( [in]int32_t in ); 
	ER	putInt64( [in]int64_t in ); 
	ER	putInt128( [in]int128_t in ); 
  
	ER	getInt8( [out]int8_t *out );
	ER	getInt16( [out]int16_t *out );
	ER	getInt32( [out]int32_t *out );
	ER	getInt64( [out]int64_t *out );
	ER	getInt128( [out]int128_t *out );

	/* ̵��������� (�侩) */
	ER	putUInt8( [in]uint8_t in ); 
	ER	putUInt16( [in]uint16_t in ); 
	ER	putUInt32( [in]uint32_t in ); 
	ER	putUInt64( [in]uint64_t in ); 
	ER	putUInt128( [in]uint128_t in ); 
  
	ER	getUInt8( [out]uint8_t *out );
	ER	getUInt16( [out]uint16_t *out );
	ER	getUInt32( [out]uint32_t *out );
	ER	getUInt64( [out]uint64_t *out );
	ER	getUInt128( [out]uint128_t *out );

	/* ʸ�����ʿ侩��8bit�� */
	ER	putChar( [in]char_t in ); 
	ER	getChar( [out]char_t *out ); 

	/* ��ư������ */
	ER	putFloat32( [in]float32_t in );
	ER	putDouble64( [in]double64_t in );
	ER	getFloat32( [out]float32_t *out );
	ER	getDouble64( [out]double64_t *out );


	/* ��侩�η�(ͭ���) */
	ER	putSChar( [in]schar_t in );
	ER	putShort( [in]short_t in ); 
	ER	putInt( [in]int_t in ); 
	ER	putLong( [in]long_t in ); 

	ER	getSChar( [out]schar_t *out ); 
	ER	getShort( [out]short_t *out ); 
	ER	getInt( [out]int_t *out ); 
	ER	getLong( [out]long_t *out ); 


	/* ��侩�η�(̵���) */
	ER	putUChar( [in]uchar_t in ); 
	ER	putUShort( [in]ushort_t in ); 
	ER	putUInt( [in]uint_t in ); 
	ER	putULong( [in]ulong_t in ); 

	ER	getUChar( [out]unsigned char *out ); 
	ER	getUShort( [out]ushort_t *out ); 
	ER	getUInt( [out]uint_t *out ); 
	ER	getULong( [out]ulong_t *out ); 

	ER	putIntptr( [in]const intptr_t ptr );
	ER	getIntptr( [out]intptr_t *ptr );
};

celltype tTDR {
	call	sChannel	cChannel;
	[inline]
		entry	sTDR	eTDR;

	var {
		TMO	tmo = C_EXP( "TMO_FEVR" );
	};
	require tSysLog.eSysLog;
};

celltype tNBOTDR {
	call	sChannel	cChannel;
	[inline]
		entry	sTDR	eTDR;

	var {
		TMO	tmo = C_EXP( "TMO_FEVR" );
	};
	require tSysLog.eSysLog;
};
