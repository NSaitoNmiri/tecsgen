/* composite ��Υ��������Υƥ��ȥ����� */
/* composite �Υ��������ˤϡ�����¾�˥�졼��������(composite_alloc2)������ե�������(composite_alloc3)������ */

import_C( "cygwin_tecs.h" );
import( "cygwin_kernel.cdl" );

/*
  1) Composite call, entry �� signature �� send/receive �������硢���������ƤӸ��ʳ��������ѡˤ���������
  2) CompositeCelltypeJoin ����������ݤ� port �� send/receive ����ľ����������˸ƤӸ��� export ������������

  080307ʸˡ�ξ��μ��������
  ����ʸˡ�Ǥ� allocator ����Ҥ���Ĺ�ʾ嵭�������Ф�̷�������å����������
  composite ����� allocator ��������ɬ�פ�����Ρ�
  (�ष����ʤ��ۤ����褤�ΤǤϤʤ���)
  1) composite_statement_specifier_list ���ߤ��� bnf.y.rb
     => ����֤���ɬ�פ���
  2) Composite call, entry �� signature �� send/receive �������硢���������ƤӸ��ʳ��������ѡˤ���������
  3) allocator �� => �ξ�� CompositecelltypeJoin ������
  
 */

signature sAlloc {
	ER  alloc( [in]int32_t size, [out]void **p );
	ER  dealloc( [in]const void *p );
};

signature sAllocTMO {
	ER  alloc( [in]int32_t size, [out]void *p, [in]TMO tmo );
	ER  dealloc( [in]const void *p );
};

celltype tAlloc {
	entry sAlloc eA;
	attr {
		int32_t  size = 8192;
	};
	var {
		[size_is(size)]
			int8_t  *buffer;
	};
};

signature sSendRecv {
	/* ���δؿ�̾�� send, receive ��ȤäƤ��ޤ��� allocator ����Ǥ��ʤ� */
	ER snd( [send(sAlloc),size_is(sz)]int8_t *buf, [in]int32_t  sz );
	ER rcv( [receive(sAlloc),size_is(*sz)]int8_t **buf, [out]int32_t  *sz );
};

celltype tTestComponent {
	entry  sSendRecv eS;
	call   sSendRecv cS;
};

celltype tTestServ {
	entry  sSendRecv eS;
};

celltype tTestClient {
	call   sSendRecv cS;
	entry  sTaskBody eBody;
};

composite tComp {
	entry sSendRecv eSe;
	call  sSendRecv cS;

	cell tTestComponent InComp{
		cS => composite.cS;
	};
	composite.eSe => InComp.eS;
};

/*
 *
 * +-------+   +------+    +----------+    +-------------+
 * |  Task | --|> Top |----|>  Middle |----|>   Bottom   |
 * +-------+   +------+  | +----------+  | +-------------+
 *                       |               |
 *                       +-------+-------+
 *                               |
 *                          +-----------+
 *                          |    V      |
 *                          |   Alloc   |
 *                          +-----------+
 */

cell tAlloc alloc {
};

[allocator(
	eS.snd.buf=alloc.eA,
	eS.rcv.buf=alloc.eA
	)]
cell tTestServ Bottom{
};

[allocator(
	eS.snd.buf=alloc.eA,
	eS.rcv.buf=alloc.eA
	)]
cell tTestComponent Middle{
	cS = Bottom.eS;
};

cell tTestClient Top {
	cS = Middle.eS;
};

[allocator(
	eSe.snd.buf=alloc.eA,
	eSe.rcv.buf=alloc.eA
	)]
cell tComp Middle2{
	cS = Bottom.eS;
};

cell tTestClient Top2 {
	cS = Middle2.eSe;
};

cell tTask Task1 {
	cBody = Top.eBody;
	priority = 1;
	stackSize = 4096;
	taskAttribute = C_EXP("TA_ACT");
};

cell tTask Task2 {
	cBody = Top2.eBody;
	priority = 1;
	stackSize = 4096;
	taskAttribute = C_EXP("TA_ACT");
};

/*
 * tCompRec: tComp ��Ƶ�Ū�� composite �ˤ������
 */
composite tCompRec {
	entry sSendRecv eSx;
	call  sSendRecv cS;
	
	cell tComp Comp {
		cS => composite.cS;
	};
	composite.eSx => Comp.eSe;
};

[allocator(
	eSx.snd.buf=alloc.eA,
	eSx.rcv.buf=alloc.eA
	)]
cell tCompRec CompRec {
	cS = Bottom.eS;
};


/*
 * �����ǥ��������˷�礷�Ƥ���ʥ�졼���Ƥ��ʤ���
 * �����ˤϷ��ϽФƤ��ʤ�
 *
 *   +----------------------------------------------+
 *   |  tTriple                                     |
 *   | +------+    +----------+    +-------------+  |
 *  -+-|> Top |----|>  Middle |----|>   Bottom   |  |
 *   | +------+  | +----------+  | +-------------+  |
 *   |           |               |                  |
 *   |           +-------+-------+                  |
 *   |                   |                          |
 *   |              +-----------+                   |
 *   |              |    V      |                   |
 *   |              |   Alloc   |                   |
 *   |              +-----------+                   |
 *   +----------------------------------------------+
 */
composite tTriple {
	entry sTaskBody eTaskBody;

	cell tAlloc Alloc {};

	[allocator(
			   eS.snd.buf=Alloc.eA,
			   eS.rcv.buf=Alloc.eA
			   )]
	cell tTestServ Bottom{
	};

	[allocator(
			   eS.snd.buf=Alloc.eA,
			   eS.rcv.buf=Alloc.eA
			   )]
	cell tTestComponent Middle{
		cS = Bottom.eS;
	};
	cell tTestClient    TopB{
		cS = Middle.eS;
	};
	composite.eTaskBody => TopB.eBody;
};

cell tTriple Triple {
};

cell tTask Task3 {
	cBody = Triple.eTaskBody;
	priority = 1;
	stackSize = 4096;
	taskAttribute = C_EXP("TA_ACT");
};


/*
 * tTriple2: tTrple �� Middle �� composite �ˤ������
 */
composite tTriple2 {
	entry sTaskBody eTaskBody;

	cell tAlloc Alloc {};

	[allocator(
			   eS.snd.buf=Alloc.eA,
			   eS.rcv.buf=Alloc.eA
			   )]
	cell tTestServ Bottom{
	};

	[allocator(
			   eSx.snd.buf=Alloc.eA,
			   eSx.rcv.buf=Alloc.eA
			   )]
	cell tCompRec Middle{
		cS = Bottom.eS;
	};
	cell tTestClient    Top{
		cS = Middle.eSx;
	};
	composite.eTaskBody => Top.eBody;
};

cell tTriple2 Triple2 {
};

cell tTask Task4 {
	cBody = Triple2.eTaskBody;
	priority = 1;
	stackSize = 4096;
	taskAttribute = C_EXP("TA_ACT");
};

