/* composite ��Υ��������Υƥ��ȥ����� */
/* composite �Υ��������ˤϡ�����¾�˥�졼��������(composite_alloc2)������ե�������(composite_alloc3)������ */

import_C( "cygwin_tecs.h" );
import( "cygwin_kernel.cdl" );

/*
  1) Composite call, entry �� signature �� send/receive �������硢���������ƤӸ��ʳ��������ѡˤ���������
  2) CompositeCelltypeJoin ����������ݤ� port �� send/receive ����ľ����������˸ƤӸ��� export ������������

  080307ʸˡ�ξ��μ��������
  ����ʸˡ�Ǥ� allocator ����Ҥ���Ĺ�ʾ嵭�������Ф�̷�������å����������
  composite ����� allocator ��������ɬ�פ�����Ρ�
  (�ष����ʤ��ۤ����褤�ΤǤϤʤ���)
  1) composite_statement_specifier_list ���ߤ��� bnf.y.rb
     => ����֤���ɬ�פ���
  2) Composite call, entry �� signature �� send/receive �������硢���������ƤӸ��ʳ��������ѡˤ���������
  3) allocator �� => �ξ�� CompositecelltypeJoin ������
  
 */

signature sAlloc {
	ER  alloc( [in]int32_t size, [out]void **p );
	ER  dealloc( [in]const void *p );
};

signature sAllocTMO {
	ER  alloc( [in]int32_t size, [out]void *p, [in]TMO tmo );
	ER  dealloc( [in]const void *p );
};

celltype tAlloc {
	entry sAlloc eA;
	attr {
		int32_t  size = 8192;
	};
	var {
		[size_is(size)]
			int8_t  *buffer;
	};
};

cell tAlloc alloc {
};

signature sSendRecv {
	/* ���δؿ�̾�� send, receive ��ȤäƤ��ޤ��� allocator ����Ǥ��ʤ� */
	ER snd( [send(sAlloc),size_is(sz)]int8_t *buf, [in]int32_t  sz );
	ER rcv( [receive(sAlloc),size_is(*sz)]int8_t **buf, [out]int32_t  *sz );
};

celltype tTestComponent {
	entry  sSendRecv eS;
	call   sSendRecv cS;
};

celltype tTestServ {
	entry  sSendRecv eS;
};

[allocator(
	eS.snd.buf=alloc.eA,
	eS.rcv.buf=alloc.eA
	)]
cell tTestServ TestServ{
};

[allocator(
	eS.snd.buf=alloc.eA,
	eS.rcv.buf=alloc.eA
	)]
cell tTestComponent comp{
	cS = TestServ.eS;
};

celltype tTestClient {
	call   sSendRecv cS;
	entry  sTaskBody eBody;
};

cell tTestClient Client1 {
	cS = comp.eS;
};

composite tComp {
	entry sSendRecv eSe;
	call  sSendRecv cS;

	cell tTestComponent comp{
		cS => composite.cS;
	};
	composite.eSe => comp.eS;
};

[allocator(
	eSe.snd.buf=alloc.eA,
	eSe.rcv.buf=alloc.eA
	)]
cell tComp Comp2{
	cS = TestServ.eS;
};

cell tTestClient Client2 {
	cS = Comp2.eSe;
};

cell tTask Task1 {
	cBody = Client1.eBody;
	priority = 1;
	stackSize = 4096;
	taskAttribute = C_EXP("TA_ACT");
};

cell tTask Task2 {
	cBody = Client2.eBody;
	priority = 1;
	stackSize = 4096;
	taskAttribute = C_EXP("TA_ACT");
};
