signature sSig1 {
  int32_t func1( [in]int32_t arg );
};


celltype tCell1 {
   call sSig1 cCall;
};

celltype tOnlyProtoCell2 {
   entry sSig1 eEnt;
};


cell tOnlyProtoCell2 cell2 ;       /* �ץ�ȥ���������Τߡ����Τ�̵�� */
cell tCell1 cellx;                 /* �ץ�ȥ���������Τߡ����Ȥ���ʤ� */

cell tCell1 cell1 {
   cCall = cell2.eEnt;
};

/* cell2 �ϥץ�ȥ���������Τߤǡ�����������ʤ�
cell tOnlyProtoCell2 cell2 {
};
 */