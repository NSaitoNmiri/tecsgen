typedef struct t_in4_ifaddr_ {
	uint32_t addr; /* IPv4 ���ɥ쥹 */
	uint32_t mask; /* ���֥ͥåȥޥ��� */
} T_IN4_IFADDR_;

signature sIfetherv4 {
	void func( void );
};

[singleton]
celltype tIfetherv4 {
	attr {
		T_IN4_IFADDR_ ether_ifnet_a = {0,0};   // ����ʤ�
	};
	var{
		T_IN4_IFADDR_ ether_ifnet_v = {0,0};   // typedef ���줿�����б��Ǥ��Ƥ��ʤ�. Ruby �㳰
	};
	[inline]entry sIfetherv4 eIfetherv4;
};

cell tIfetherv4 Ifetherv4 {
	
};
