/*
 *  ���ꥢ�륤�󥿥ե������ɥ饤�Ф�ư�������ѤΤ�������
 *
 *  �ʲ�������ϡ��ӥå���������¤�Ȥä��Ѥ��롥
 */
const unsigned int IOCTL_NULL	=0;		/* ����ʤ� */
const unsigned int IOCTL_ECHO	=0x0001;		/* ��������ʸ���򥨥����Хå� */
const unsigned int IOCTL_CRLF	=0x0010;		/* LF �������������� CR ���ղ� */
const unsigned int IOCTL_FCSND	=0x0100;		/* �������Ф��ƥե������Ԥ� */
const unsigned int IOCTL_FCANY	=0x0200;		/* �ɤΤ褦��ʸ���Ǥ������Ƴ� */
const unsigned int IOCTL_FCRCV	=0x0400;		/* �������Ф��ƥե������Ԥ� */

/*
 *  ������μ��̤����
 *
 *  LOG_TYPE_CYC��LOG_TYPE_ASSERT �ʳ��ϡ��ǥХå��󥰥��󥿥ե�������
 *  �ͤȹ��פ��Ƥ��롥
 */
const unsigned int LOG_TYPE_INH	=	0x01;	/* ����ߥϥ�ɥ� */
const unsigned int LOG_TYPE_ISR	=	0x02;	/* ����ߥ����ӥ��롼���� */
const unsigned int LOG_TYPE_CYC	=	0x03;	/* �����ϥ�ɥ� */
const unsigned int LOG_TYPE_EXC	=	0x04;	/* CPU�㳰�ϥ�ɥ� */
const unsigned int LOG_TYPE_TEX	=	0x05;	/* �������㳰�����롼���� */
const unsigned int LOG_TYPE_TSKSTAT =	0x06;	/* �����������Ѳ� */
const unsigned int LOG_TYPE_DSP	=	0x07;	/* �ǥ����ѥå��� */
const unsigned int LOG_TYPE_SVC	=	0x08;	/* �����ӥ������� */
const unsigned int LOG_TYPE_COMMENT =	0x09;	/* ������ */
const unsigned int LOG_TYPE_ASSERT =	0x0a;	/* �����������μ��� */

const unsigned int LOG_ENTER	=	0x00;	/* ���������� */
const unsigned int LOG_LEAVE	=	0x80;	/* �и�����λ */

/*
 *  ������ν����٤����
 */
const unsigned int LOG_EMERG	=0;		/* ����åȥ�������ͤ��륨�顼 */
const unsigned int LOG_ALERT	=1;
const unsigned int LOG_CRIT	=2;
const unsigned int LOG_ERROR	=3;		/* �����ƥ२�顼 */
const unsigned int LOG_WARNING	=4;		/* �ٹ��å����� */
const unsigned int LOG_NOTICE	=5;
const unsigned int LOG_INFO	=6;
const unsigned int LOG_DEBUG	=7;		/* �ǥХå��ѥ�å����� */


const int TMAX_LOGINFO	= 6;
/* #define TMAX_LOGINFO 6 */

 const int NULL = 0;
 const int FALSE = 0;
 const int32 SERIAL_BUFSZ = 256;
 const int32 SERIAL_RCV_SEM1 = 1;
 const int32 SERIAL_SND_SEM1 = 2;
 const int32 SERIAL_RCV_SEM2 = 3;
 const int32 SERIAL_SND_SEM2 = 4;

 /*��
 	����� 
 	       �������ؿ��Ȥ���
 	       Factory�ǻ��ꤹ��
 	       ITRON�Ǥ���ŪAPI�ǽ�����ϥ�ɥ�˻��ꤹ��
 	       

 */


 /*
 	LogOutput����Ȥ��ƤϽ������ɬ�פʤ�
 	sio_initialize()��SerialIOPort����ν�����Ǥ���
 	����ȥ���֥�å��ν�����ϡ����ꥢ��ݡ��ȥ����°�����ѿ�
 	�ν�����Ǽ¸�����
 	�ݡ��Ȥν�����ϥ������³����ꤷ���Ȥ�����ޤ�

 	����Ū��(���뤤�����Ū��)�����Ϥξ��֤λ��ȤϽ��褿�Ȥ��Ƥ⡢
 	���ꥢ��ݡ�����ͭ�ξ��֤ι��ܤλ��Ȥϡ�����Ū�ʥ����Ϥξ���
 	���Ȥ���ϡ�ľ�ܻ���Ǥ��ʤ��ΤǤ�̵����?
 */


 /****/

 /* for SH3 */
 typedef signed   int32	INT;
 typedef signed   int32	SYSTIM;
 typedef signed   int32	VP_INT;
 typedef unsigned int32	UINT;
 typedef unsigned int32	UW;
 typedef unsigned int8	UB;

 /* for uITRON4.0 */

 typedef INT		ER;
 typedef INT		ID;
 typedef INT		ER_UINT;
 typedef bool		BOOL;


 /* for serial */
 /*
  *  ���ꥢ��ݡ��ȴ����֥�å�
  */

 typedef struct serial_port_initialization_block {
 	ID	rcv_semid;	/* �����Хåե������ѥ��ޥե���ID */
 	ID	snd_semid;	/* �����Хåե������ѥ��ޥե���ID */
 } SPINIB;

 typedef struct serial_port_control_block {
 	BOOL	openflag;	/* �����ץ�Ѥߥե饰 */
 	UINT	ioctl;		/* ư������������� */

 	UINT	rcv_read_ptr;	/* �����Хåե��ɽФ��ݥ��� */
 	UINT	rcv_write_ptr;	/* �����Хåե�����ߥݥ��� */
 	UINT	rcv_count;	/* �����Хåե����ʸ���� */
 	char	rcv_fc_chr;	/* ����٤� START/STOP */
 	BOOL	rcv_stopped;	/* STOP �����ä����֤��� */

 	UINT	snd_read_ptr;	/* �����Хåե��ɽФ��ݥ��� */
 	UINT	snd_write_ptr;	/* �����Хåե�����ߥݥ��� */
 	UINT	snd_count;	/* �����Хåե����ʸ���� */
 	BOOL	snd_stopped;	/* STOP �������ä����֤��� */

 	char	rcv_buffer[SERIAL_BUFSZ];	/* �����Хåե� */
 	char	snd_buffer[SERIAL_BUFSZ];	/* �����Хåե� */
 } SPCB;

 /*
  *  ���ꥢ�륤�󥿥ե������ɥ饤�Ф��Ѥ���ѥ��å�
  */
 typedef struct {
 	UINT	reacnt;		/* �����Хåե����ʸ���� */
 	UINT	wricnt;		/* �����Хåե����ʸ���� */
 } T_SERIAL_RPOR;

 const int32 SIO_ERDY_SND = 0;   /* oyama */
 const int32 SIO_ERDY_RCV = 1;

 /*
  *  ���ꥢ��I/O�ݡ��Ƚ�����֥�å�
  */
 typedef struct sio_port_initialization_block {
     UW reg_base;    /* �쥸�����Υ١������ɥ쥹 */
     UB lcr_val;     /* �⡼�ɥ쥸������������   */
     UB dlm_val;     /* �ܡ��졼�Ⱦ�̤�������   */
     UB dll_val;     /* �ܡ��졼�Ȳ��̤�������   */
     UW pinter_val;  /* ����ߵ��ĥӥå�   */    
 } SIOPINIB;

 /*
  *  ���ꥢ��I/O�ݡ��ȴ����֥�å�
  */
 typedef struct {
     VP_INT  exinf;		/* ��ĥ���� */
     BOOL    openflag;		/* �����ץ�Ѥߥե饰 */
     BOOL    sendflag;		/* ��������ߥ��͡��֥�ե饰 */
     BOOL    getready;		/* ʸ��������������� */
     BOOL    putready;		/* ʸ���������Ǥ������ */
 } SIOPCB;

typedef struct {
	UINT	logtype;		/* ������μ��� */
	SYSTIM	logtim;			/* ������ */
	VP_INT	loginfo[TMAX_LOGINFO];	/* ����¾�Υ����� */
} SYSLOG;


signature sLog {
	  void log(void);	
};

signature sSysLog {
	  ER vwri_log( [in] UINT prio,  [in] SYSLOG *p_log);
	  ER_UINT vrea_log( [out] SYSLOG *p_log);
	  ER vmsk_log( [in] UINT logmask,  [in] UINT lowmask);

	  ER opn_port( void ); /* �ݡ��ȤΥ����ץ� */
	  ER cls_port( void ); /* �ݡ��ȤΥ����� */
};

const int TCNT_SYSLOG_BUFFER = 32;

signature sFormattedOutput {
	  void syslog_output( void );
	  void syslog_print( [in] SYSLOG *p_log );
	  void syslog_printf( [in,string] char *format, [in,size_is(expr)] VP_INT *args, [in] int expr);

 	  ER opn_port( void ); /* �ݡ��ȤΥ����ץ� */
 	  ER cls_port( void ); /* �ݡ��ȤΥ����� */
 	  ER_UINT wri_dat( [in , size_is(len)] char *buf,  [in] UINT len); /* ʸ������
 	  �� */
 	  ER_UINT rea_dat( [out , size_is(len)] char *buf,  [in] UINT len); /* ʸ����
 	  ���� */
 	  ER ctl_por( [in] UINT ioctl); /* �ݡ��Ȥ����� */
};

signature sPort {
 	  ER opn_port( void ); /* �ݡ��ȤΥ����ץ� */
 	  ER cls_port( void ); /* �ݡ��ȤΥ����� */
 	  ER_UINT wri_dat( [in , size_is(len)] char *buf,  [in] UINT len); /* ʸ������
 	  �� */
 	  ER_UINT rea_dat( [out , size_is(len)] char *buf,  [in] UINT len); /* ʸ����
 	  ���� */
 	  ER ctl_por( [in] UINT ioctl); /* �ݡ��Ȥ����� */

};


signature sSerialPortCallBack {
 	  void ierdy_snd( [in] VP_INT exinf);/* ���ꥢ��ݡ��Ȥ����������ǽ������Хå� */
 	  void ierdy_rcv( [in] VP_INT exinf); /* ���ꥢ��ݡ��Ȥ���μ������Υ�����Хå� */
};

signature sSIOPort {
 	  void opn_por( [in] ID id , [in] VP_INT exinf);
 	  void cls_por( [in] ID id);
 	  BOOL snd_chr( [in] char c);
 	  INT  rcv_chr( void );
 	  void ena_cbr( [in] UINT cbrtn);
 	  void dis_cbr( [in] UINT cbrtn);
 	  void init_for_banner(void);

 	  /* ������ϥ�ɥ� */
 	  void initialize(void);
 	  /* ����ߥϥ�ɥ� */
 	  void interrupt(void);
};

[singleton] 
celltype tLog {
	entry sLog eLog;
	call  sFormattedOutput cFormattedOutput;
};

[singleton] 
celltype tSysLog {
	entry sSysLog eSysLog;
	call  sFormattedOutput cFormattedOutput;

	  var {
	  /*
	   *  ���Ϥ��٤�������ν����١ʥӥåȥޥåס�
	    */
	    UINT	syslog_logmask;			/* ���Хåե��˵�Ͽ���٤������� */
	    UINT	syslog_lowmask;			/* ���٥���Ϥ��٤������� */
	  /*
	   *  ���Хåե��Ȥ���˥����������뤿��Υݥ���
	    */
	     SYSLOG	syslog_buffer[TCNT_SYSLOG_BUFFER];	/* ���Хåե� */
	     UINT	syslog_count;			/* ���Хåե���Υ��ο� */
	     UINT	syslog_head;			/* ��Ƭ�Υ��γ�Ǽ���� */
	     UINT	syslog_tail;			/* ���Υ��γ�Ǽ���� */
	     UINT	syslog_lost;			/* ����줿���ο� */
	  };

 /*
 �ʲ��δؿ��ϼ���ȼ����ɲä���

	 factory( INIT_HANDLER ,      TA_HLG, 0, tSysLog_initialize );
 	 factory( INTERRUPT_HANDLER , TA_HLG, INHNO_SIO, tSysLog_interrupt );*/

};

celltype tFormattedOutput {
	entry  sFormattedOutput eFormattedOutput;
	call   sPort cPort;
	call   sSysLog cSysLog;
};

celltype tLowOutputSIO {
	entry sPort ePort;
	call  sSIOPort cSIOPort;
};

celltype tSerialPort {
	entry sPort ePort;
	entry sSerialPortCallBack eSerialPortCallBack;
	call  sSIOPort cSIOPort;

	var {
		SPCB spcb;
	};
};

celltype tSIOPortLinux {
	entry sSIOPort eSIOPort;
	call sSerialPortCallBack cSerialPortCallBack;

	var {
		SIOPCB siopcb;
	};
};

celltype tSIOPortST16C2550 {
	entry sSIOPort eSerialIOPort[2];
	call sSerialPortCallBack eSerialPortCallBack;

	var {
		SIOPCB siopcb;
	};
};

 /* �ץ�ȥ�������� */
cell tSerialPort SerialPort;

cell tSIOPortLinux SIOPortLinux {
	cSerialPortCallBack = SerialPort.eSerialPortCallBack;

/*      siopcb = { {FALSE,FALSE,FALSE,FALSE},
                 {FALSE,FALSE,FALSE,FALSE}
		 };      060830 */
/*
      siopinib = { {ST16C_CHB, LCR_VAL, DLM_VAL, DLL_VAL, PINTER_PINT7E},
 		   {ST16C_CHA, LCR_VAL, DLM_VAL, DLL_VAL, PINTER_PINT6E}
 		   };
*/
};

cell tSerialPort SerialPort {
	cSIOPort = SIOPortLinux.eSIOPort;
      	spcb = { FALSE , 0 , NULL , NULL, 0 , '\0' , FALSE };
      /*spinib = { SERIAL_RCV_SEM1, SERIAL_SND_SEM1 };  060830 */
};



/* cell tSIOPortST16C2550 SIOPortST16C2550;
*/
cell tLowOutputSIO LowOutputSIO {
	cSIOPort = SIOPortLinux.eSIOPort;
};

/* 
cell tLowOutputSTUB LowOutputSTUB{
	cPort = SIOPortLinux.eSIOPort;
};
*/
cell tFormattedOutput FormattedOutputSysLog {
	cPort = LowOutputSIO.ePort;
};

cell tFormattedOutput FormattedOutput {
	cPort = SerialPort.ePort;
};

cell tSysLog SysLog {
	cFormattedOutput = FormattedOutputSysLog.eFormattedOutput;
};

cell tLog Log {
	  cFormattedOutput = FormattedOutput.eFormattedOutput;
};



