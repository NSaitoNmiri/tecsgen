import_C( "tecs.h" );
/* typedef int32_t ER; */

const int32_t  const_int = 32;

signature sSig {
	/* ER func( [in]int32_t in, [out]int32_t *out ); */
	int32_t func( [in]int32_t in, [out]int32_t *out );
};

celltype tCt {
	entry  sSig eEnt;
	attr {
		int32_t  a = 20;
	};
	var {
		int32_t  v = 31;
	};
};


cell tCt C0 {};
cell tCt C1 {};


celltype tCt2 {
	call sSig cCall0;
	call sSig cCall1;

	attr {
		int32_t  a = 20;
	};
	var {
		int32_t  v = 31;
	};
 
};

cell tCt2 ct2 {
  cCall0 = C0.eEnt;
  cCall1 = C1.eEnt;
};


celltype tOmit{
	attr {
		[omit]int32_t  a;
	};
	factory{
		write( "tecsgen.cfg", "tOmit cb=$cb$ id=$id$ idx=$idx$ ID=$ID$" );
	};
};

cell tOmit om1
{
	a = -100;
};

[idx_is_id]
celltype tIdx_is_id {
	entry sSig eEnt;
	attr {
		int32_t  a_init = 10;
		int32_t  b_init = -20;
		int32_t  c_init;
	};
	var {
		int32_t  a = a_init;
		int32_t  b = b_init + 1;
		int32_t  c = c_init * 2;
	};
	factory{
		write( "tecsgen.cfg", "tIdx_is_id cb=$cb$ id=$id$ idx=$idx$ ID=$ID$" );
	};
};

cell  tIdx_is_id cell_idx_is_id1 {
	a_init = 100;
	c_init = -40;
};

cell  tIdx_is_id cell_idx_is_id2 {
	b_init = -200;
	c_init = -50;
};

cell  tIdx_is_id cell_idx_is_id3 {
	c_init = 1000;
};

[singleton,idx_is_id]
celltype tSingle_idx_is_id {
	factory {
		write( "tecsgen.cfg", "tSingle_idx_is_id cb=$cb$ id=$id$ idx=$idx$ ID=$ID$" );
	};
};

cell tSingle_idx_is_id cell_single {
};

celltype tVarInitByAttr {
	attr {
		int32_t   a0 = 10 + const_int;
		int32_t   a1;
	};
	var {
		int32_t   v0 = a0;
		int32_t   v1 = a1 + const_int;
	};
	entry sSig eEnt;
};

cell tVarInitByAttr Cell1 {
	a1 = 20;
};

cell tVarInitByAttr Cell2 {
	a0 = 101;
	a1 = 100;
};

[singleton]
celltype tSingle {
	entry sSig eSig;
	call  sSig cCall[];
	attr {
		int32_t a = 33;
	};
	var {
		int32_t b = 44;
	};
};

cell tSingle Single {
	cCall[] = Cell1.eEnt;
	cCall[] = Cell2.eEnt;
};

/* 2.  size_is �դ��� var ����������������뤫�Υƥ��� */

/* 2.1 singleton �ξ�� */
/* 2.1.1 CB, INIB �Ȥ�ˤʤ�(������ INIB �� buf �Ͻ��� */
[singleton]
celltype tSCt_no_CB_no_INIB {
	var {
		[size_is(1)]
			int8_t    *buf;
	};
};
cell tSCt_no_CB_no_INIB SCt_no_CB_no_INIB {};

/* 2.1.2 CB ����, INIB �ʤ�(������ INIB �� buf �Ͻ��� */
[singleton]
celltype tSCt_a_CB_no_INIB {
	var {
		int32_t    a = 5;
		[size_is(1)]
			int8_t    *buf;
	};
};
cell tSCt_a_CB_no_INIB SCt_a_CB_no_INIB {};

/* 2.1.3 CB �ʤ�, INIB ���� */
[singleton]
celltype tSCt_no_CB_a_INIB {
	attr {
		int32_t    size = 6;
	};
	var {
		[size_is(size)]
			int8_t    *buf;
	};
};
cell tSCt_no_CB_a_INIB SCt_no_CB_a_INIB {};

/* 2.1.3 CB, INIB �Ȥ�ˤ��� */
[singleton]
celltype tSCt_a_CB_a_INIB {
	attr {
		int32_t    size = 6;
	};
	var {
		int32_t    a = 9;
		[size_is(size)]int8_t    *buf;
	};
};
cell tSCt_a_CB_a_INIB SCt_a_CB_a_INIB {};

/* 2.2 �� singleton �ξ�� */
/* 2.2.1 CB, INIB �Ȥ�ˤʤ�(������ INIB �� buf �Ͻ��� */
celltype tCt_no_CB_no_INIB {
	var {
		[size_is(1)]int8_t    *buf;
	};
};
cell tCt_no_CB_no_INIB Ct_no_CB_no_INIB {};

/* 2.2.2 CB ����, INIB �ʤ�(������ INIB �� buf �Ͻ��� */
celltype tCt_a_CB_no_INIB {
	var {
		int32_t    a = 5;
		[size_is(1)]int8_t    *buf;
	};
};
cell tCt_a_CB_no_INIB Ct_a_CB_no_INIB {};

/* 2.2.3 CB �ʤ�, INIB ���� */
celltype tCt_no_CB_a_INIB {
	attr {
		int32_t    size = 6;
	};
	var {
		[size_is(size)]int8_t    *buf;
	};
};
cell tCt_no_CB_a_INIB Ct_no_CB_a_INIB {};

/* 2.2.3 CB, INIB �Ȥ�ˤ��� */
celltype tCt_a_CB_a_INIB {
	attr {
		int32_t    size = 6;
	};
	var {
		int32_t    a = 9;
		[size_is(size)]int8_t    *buf;
	};
};
cell tCt_a_CB_a_INIB Ct_a_CB_a_INIB {};

/* 2.3.1 CB, INIB �Ȥ�ˤʤ�(������ INIB �� buf �Ͻ���)��buf �˽����ͭ */
celltype tCt_no_CB_no_INIB_init {
	var {
		[size_is(2)]int8_t    *buf = { 99, -99 };
	};
};
cell tCt_no_CB_no_INIB_init Ct_no_CB_no_INIB_init {};

[singleton]
celltype tMain{
	call sSig cSig[];
/*
	attr {
		int32_t  a;
	};
*/
};

cell tMain MainCell {
	cSig[] = Single.eSig;
	cSig[] = C0.eEnt;
/*	cSig[2] = Cell1.eEnt;
	cSig[3] = Cell2.eEnt; */

/* */
};

