import_C( "cygwin_tecs.h" );

////////////////////////////////

typedef struct tagSt {
	int32_t		m;
} ST;

signature sTest {
	void		test( [in]int_t input );
	int32_t		test2( [in]int_t input,				[out]int32_t *ret );
	int32_t		test3( [in]const char_t *input,		[out]int32_t *ret );
	int32_t		test4( [in,string(len)]const char_t *input, [in]int32_t len );
	int32_t		test5( [in]const ST *input );
};

celltype tTECSTest {
	entry sTest eTest;
};

cell tTECSTest TECSTest {
};

// generate( RTMBridgePlugin, sTest, "\\'" );
generate( RTMBridgePlugin, sTest, "\'" );

cell tRTMsTestBridge RTMTest {
	cTECS = TECSTest.eTest;
};

// #833 $B$N%F%9%H(B $B%W%i%0%$%s@8@.$5$l$?(B cdl $B$NCf$+$i(B import( <....cdl> ); $B$5$l$F$$$k$b$N$N%;%k%?%$%W%3!<%I$r@8@.$7$F$7$^$&(B
cell tA A {
};
