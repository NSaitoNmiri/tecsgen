typedef int32_t ER;

signature sSig {
  ER func1( [in]int32_t arg1 );
  ER func2( [in]int32_t arg1 );
};

celltype tCt {
  entry sSig c;
  attr {
    int32_t a;
    int32_t ab;
    char_t *s;
    bool_t  boo = true;
  };
  var {
    int32_t b;
  };
  FACTORY {
    write( "tecs.cfg", "ATR_INI(TA_HLG, 0, tSyslog_initialize);" );
  };

  factory {
    write( "tecs.cfg", "ATR_INI(TA_HLG, 0, tSyslog_initialize);" );
    write( "tecs.cfg", "a = %d;, %d;, %s; ", a, ab, s );
    write( "tecs.cfg", "a = %d;, %d;, %s;", a, ab, s );

    write( "tecs.cfg", "a = %d;, %d;, %s; %d", a, ab, s, boo );  /* boo �� %d ���б� */
    write( "tecs.cfg", "a = %d;, %d;, %s; %d %d %s", a, ab, s );  /* %s ��¿���� */

  };
};

cell tCt ce {
  a = 0;
  ab = 99;
  s = "abc";
};
