import_C( "tecs.h" );

signature sSig{
  void func( void );
};

/*** 1.ñ�쥻���Ŭ�� ***/
// ñ�쥻���Ŭ�� (VMT ���׺�Ŭ����������ȥ����׺�Ŭ����ޤ�)
// ����¦�Υ��뤬��Ĥǡ��ݡ��Ȥ��Ĥ���

celltype tSingleCellOptimizeCaller {
  call sSig cCall;
  entry sSig eEnt;
};

celltype tSingleCellOptimizeCallee {
  entry sSig eEnt;
};

// �Ƥ�¦���� 1����
cell tSingleCellOptimizeCallee SingleCellOptimizeCallee;

cell tSingleCellOptimizeCaller SingleCellOptimizeCaller {
  cCall = SingleCellOptimizeCallee.eEnt;
};
// ����¦����
cell tSingleCellOptimizeCallee SingleCellOptimizeCallee {
};
// �Ƥ�¦���� 2����
cell tSingleCellOptimizeCaller SingleCellOptimizeCaller2 {
  cCall = SingleCellOptimizeCallee.eEnt;
};

/*** 2. VMT ���׺�Ŭ�� ***/
// ����¦�Υ��뤬��Ĥ���������������

celltype tVMTUselessOptimizeCaller {
  call sSig cCall;
  entry sSig eEnt;
};

celltype tVMTUselessOptimizeCallee {
  entry sSig eEnt[2];
  attr {
	  int32_t  attribute = 100;
  };
};

// ����¦����
cell tVMTUselessOptimizeCallee VMTUselessOptimizeCallee;

// �Ƥ�¦���� 1����
cell tVMTUselessOptimizeCaller VMTUselessOptimizeCaller {
  cCall = VMTUselessOptimizeCallee.eEnt[0];
};
// �Ƥ�¦���� 2����
cell tVMTUselessOptimizeCaller VMTUselessOptimizeCaller2 {
  cCall = VMTUselessOptimizeCallee.eEnt[1];
};
// ����¦����
cell tVMTUselessOptimizeCallee VMTUselessOptimizeCallee {
};

/*** VMT ���׺�Ŭ��&������ȥ����׺�Ŭ�� ***/
// ����¦�Υ��뤬ʣ��������ñ��Υ��륿����

celltype tSkeltonUselessOptimizeCaller {
  call sSig cCall;
  entry sSig eEnt;
};

celltype tSkeltonUselessOptimizeCallee {
  entry sSig eEnt;
  attr {
	  int32_t  attribute = 100;
  };
};

// ����¦����
cell tSkeltonUselessOptimizeCallee SkeltonUselessOptimizeCallee;
cell tSkeltonUselessOptimizeCallee SkeltonUselessOptimizeCallee2;

// �Ƥ�¦���� 1����
cell tSkeltonUselessOptimizeCaller SkeltonUselessOptimizeCaller {
  cCall = SkeltonUselessOptimizeCallee.eEnt;
};
// �Ƥ�¦���� 2����
cell tSkeltonUselessOptimizeCaller SkeltonUselessOptimizeCaller2 {
  cCall = SkeltonUselessOptimizeCallee2.eEnt;
};
// ����¦����
cell tSkeltonUselessOptimizeCallee SkeltonUselessOptimizeCallee {
};
cell tSkeltonUselessOptimizeCallee SkeltonUselessOptimizeCallee2 {
};

[singleton]
celltype tMain {
	call sSig cMain[];
};
cell tMain Main{
	cMain[0] = SingleCellOptimizeCaller.eEnt;
	cMain[1] = VMTUselessOptimizeCaller.eEnt;
    cMain[2] = SkeltonUselessOptimizeCallee.eEnt;
    cMain[3] = SkeltonUselessOptimizeCallee2.eEnt;
};

