

signature sSingleCall {
  /* int32  single( [in]int32 single );    060827   ���顼�ˤʤ�ʤ�*/
  int32  single( [in]int32 s );
};

signature sSingleEntry {
  int32  single( [in]int32 s );
};

[singleton]
celltype tSingle {
  call  sSingleCall  cCall;
  entry sSingleEntry eEntry;

  attr {

    int32  single;
  };

  var {
    int32  single_var;
  };

};

celltype tSingleCall{
  call sSingleEntry cSingleEntry;
};

celltype tSingleEntry{
  entry sSingleCall eSingleCall;
  attr{
    int32 a;
  };
};


cell tSingleEntry singleentry{
  a = 0;
};

cell tSingle single{
  cCall = singleentry.eSingleCall;
  single = 0;
};

cell tSingle single2{
  cCall = singleentry.eSingleCall;
  single = 0;
};

cell tSingleCall singlecall{
  cSingleEntry = single.eEntry;
};

composite tSingleComp {
  cell tSingle c{
    single = 10;
  };
  cSingle = c.cCall;
};

cell tSingleComp singleComp1 {
  cSingle = single.eEntry;
 };
cell tSingleComp singleComp2 {
  cSingle = single.eEntry;
};


