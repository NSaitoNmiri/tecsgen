celltype tAttr {
	attr {
		int		*a={ 1, 2 };     // �����顼�̤ʤΤǡ��ǽ����ʬ�Τߤ��Ѥ�����ˡ��ͤ����뤬���顼�Ȥ���
		[omit]
			int		b[] = { 1, 2 };  // omit ���ꤵ��Ƥ���Х��顼�ǤϤʤ�
	};
	var {
		// [size_is(*a)]		// �����㳰
		[size_is(2)]
			int8_t	*c;
	};
	factory {
		write( "tecsgen.cfg", "%s", b );
	};
};

cell tAttr Attr {
};

celltype tAttr2 {
	attr {
		int		a=10;
	};
	var {
		[size_is(a)]
			int8_t	*b;
	};
};

cell tAttr Attr2 {
};

