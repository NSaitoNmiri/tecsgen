const PRI  MAIN_PRIORITY =  5;		/* �ᥤ�󥿥�����ͥ���� */
					/* HIGH_PRIORITY ���⤯���뤳�� */
const PRI  HIGH_PRIORITY =  9;		/* ����˼¹Ԥ���륿������ͥ���� */
const PRI  MID_PRIORITY  = 10;
const PRI  LOW_PRIORITY  = 11;

/* �����ϥ�ɥ� */
[singleton]
celltype tCycMain {
  entry sMain eMain;
  call  siSystem ciSys;   /* tSampleMain �θƤӸ���̾�����Ѥ��Ƥ��� */
};

cell tCycMain cyc_main {
  ciSys = toppers_jsp.eiSystem;
};

cell tCyc cyc_hdlr {
  cHdlr = cyc_main.eMain;
  cyctim = 2000;
  cycatr = TA_HLNG;
};

/* ���֥ᥤ�󥿥��� */
[singleton]
celltype tSubMain {
  entry sMain eSubMain;
  call  sSystem cSysSub;   /* tSampleMain �θƤӸ���̾�����Ѥ��Ƥ��� */
};

cell tSubMain sub_main{
  cSysSub = toppers_jsp.eSystem;
};

cell tTask task0 {
  cMain = sub_main.eSubMain;
  exinf = 1;
  tskatr = TA_HLNG;
  itskpri = MID_PRIORITY;
};

cell tTask task1 {
  cMain = sub_main.eSubMain;
  exinf = 2;
  tskatr = TA_HLNG;
  itskpri = MID_PRIORITY;
};

cell tTask task2 {
  cMain = sub_main.eSubMain;
  exinf = 3;
  tskatr = TA_HLNG;
  itskpri = MID_PRIORITY;
};

/* �ᥤ�󥿥��� */
[singleton]
celltype tSampleMain {
  entry sMain   eMain;
  call  sTask   cTask[3];
  call  sSystem cSysMain;
  call  sCyc    cCyc;
};

cell tSampleMain sample_main {
  cTask[0]  = task0.eT;
  cTask[1]  = task1.eT;
  cTask[2]  = task2.eT;
  cSysMain  = toppers_jsp.eSystem;
  cCyc      = cyc_hdlr.eCyc;
};

cell tTask main {
  cMain = sample_main.eMain;
  tskatr = TA_HLNG | TA_ACT;
  itskpri = MAIN_PRIORITY;
};

