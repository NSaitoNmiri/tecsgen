/*
 * through �ץ饰����λ
 *
 * ��ΥХꥨ�������
 * ���������������� Plugin1, Plugin2 ��ɸ��� TracePlugin ��ľ����������롣
 *   (TracePlugin �λ�ѤǤ⤢��)
 * ��send/receive �ʥ���������
 * ��composite ���륿���פΥ���θƤӸ�
 * ���ƤӸ�����
 */
import_C( "cygwin_tecs.h" );
import( "tSysLog.cdl" );
import( "cygwin_kernel.cdl" );

struct tag { int32_t member; };
typedef int32_t INT;
typedef struct tag stTag;

signature sAlloc {
  ER    alloc( [in]int32_t sz, [out]void **ptr );
  ER    dealloc( [in]const void *ptr );
};

[singleton]
celltype tAlloc {
  entry sAlloc eA;
  var {
    int32_t  n_alloc;
    int32_t  n_dealloc;
  };
};

signature sSignature {
	ER	func1( [in]int32_t inval );
	ER	func2( [out]int32_t *outval );
	ER	func3( [in]struct tag stval );
	ER	func4( [in]stTag stval, [in]INT inval );
	ER	func5( [inout]stTag *stval, [in]INT inval );
	ER	func6( [send(sAlloc),size_is(sz)]int8_t *buf, [in]int32_t sz );
	ER	func7( [receive(sAlloc),size_is(*sz)]int8_t **buf, [out]int32_t *sz );
};

signature sSig {
	ER	func1(void );
};

signature sMain {
	ER	main( void );
};

celltype tClient {
	call	sSignature	cCall;
	call	sSignature	cCall2[2];
	entry	 sMain		eMain;
};

composite tClientComposite{
	call	sSignature	cCall;
	call	sSignature	cCall2[2];
	entry	sMain		eMain;

	cell tClient Cell {
		cCall  => composite.cCall;
		cCall2 => composite.cCall2;
	};
	composite.eMain => Cell.eMain;
};

celltype tServer {
	entry	sSignature	eEntry;
};

celltype tMain {
	call sMain cMain;
};

cell tMain Main {
	cMain = Client.eMain;
};

/*
 * ��through �λ���ˤ�ꡢplugin �ˤ����������륻��� call port �� entry port �δ֤���������
 * ��through ���������� �ץ饰����̾�����
 * ��through ����������� ���ΰ��������
 * �������ͥ졼���� through �����Ĥ��ä���硢plugin ��ƽФ� CDL ������������
 * �������ͥ졼���� through ��ޤॻ����ɤ߹�����Ȥ���ǡ��������줿 CDL ���ɤ߹�����̤Υѡ�������ѡ�
 * �����κ� typedef, signature, celltype �ϡ��ޤä���Ʊ���Ǥ���н�ʣ����Ǥ�̵�뤹��
 * ��through ��ʣ������Ǥ��������ͥ졼���ϻ��ꤵ�줿��˥������������
 * ��plugin �⥸�塼��ϡ��ƥ�ץ졼�ȥ����ɤ˴����� celltype �����ɤ��������롥
 *   (generate.rb �� gen_template_ep_fun ����������᥽�åɤ򵭽Ҥ���)
 */

cell tClientComposite Client {
//cell tClient Client {
	[ through( Plugin1, "" ),
	  through( Plugin2, "" ),
	  through( TracePlugin, "maxArrayDisplay=256" ) ]
		cCall = server.eEntry;

	[ through( Plugin1, "" ),
	  through( Plugin2, "" ),
	  through( TracePlugin, "maxArrayDisplay=64" ),
	  through( TracePlugin, "maxArrayDisplay=128" ) ]
		cCall2[0] =  server.eEntry;
	cCall2[1] =  server.eEntry; 
 };

[allocator(
		   eEntry.func6.buf=Alloc.eA,
		   eEntry.func7.buf=Alloc.eA
		   )]
cell tServer server {
};


cell tAlloc Alloc {
};

cell tSysLog SysLog {
};

cell tKernel Kernel {
};
