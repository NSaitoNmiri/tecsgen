// #833 $B$N%F%9%H(B
celltype tA {
	factory {
		write( "tecsgen.cfg", "hello!" );
	};
};
